//------------------------------------------------------------
//   Copyright 2010-2018 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------

//
// Class Description:
//
//
class apb_slave_agent_config extends uvm_object;

localparam string s_my_config_id = "apb_slave_agent_config";
localparam string s_no_config_id = "no config";
localparam string s_my_config_type_error_id = "config type error";

// UVM Factory Registration Macro
//
`uvm_object_utils(apb_slave_agent_config)

// Virtual Interface
virtual apb_slave_driver_bfm  drv_bfm;
virtual apb_slave_monitor_bfm mon_bfm;

//------------------------------------------
// Data Members
//------------------------------------------
// Is the agent active or passive
uvm_active_passive_enum active = UVM_ACTIVE;

logic[31:0] start_address[15:0];
logic[31:0] range[15:0];

int apb_index = 0;
//------------------------------------------
// Methods
//------------------------------------------
extern static function apb_slave_agent_config get_config( uvm_component c );
// Standard UVM Methods:
extern function new(string name = "apb_slave_agent_config");

//
// Task: wait_for_reset
//
// This method waits for the end of reset. 
event wait_for_reset_event;
bit   wait_for_reset_called = 0;
 
task wait_for_reset();
  if (!wait_for_reset_called) begin
    wait_for_reset_called = 1;
    mon_bfm.wait_for_reset();
    -> wait_for_reset_event;
    wait_for_reset_called = 0;
  end else begin
    @(wait_for_reset_event);
  end
endtask : wait_for_reset

endclass: apb_slave_agent_config

function apb_slave_agent_config::new(string name = "apb_slave_agent_config");
  super.new(name);
endfunction

//
// Function: get_config
//
// This method gets the my_config associated with component c. We check for
// the two kinds of error which may occur with this kind of
// operation.
//
function apb_slave_agent_config apb_slave_agent_config::get_config( uvm_component c );
  uvm_object o;
  apb_slave_agent_config t;

  if(! uvm_config_db #(uvm_object)::get(c, "", s_my_config_id, o)) begin
    c.uvm_report_error( s_no_config_id ,
                        $sformatf("no config associated with %s" ,
                                  s_my_config_id ) ,
                        UVM_NONE , `uvm_file , `uvm_line  );
    return null;
  end

  if( !$cast( t , o ) ) begin
    c.uvm_report_error( s_my_config_type_error_id ,
                        $sformatf("config %s associated with config %s is not of type my_config" ,
                                   o.sprint() , s_my_config_id ) ,
                        UVM_NONE , `uvm_file , `uvm_line );
  end

  return t;
endfunction
