//------------------------------------------------------------
//   Copyright 2010-2018 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------
package mem_ss_test_lib_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

import ahb_agent_pkg::*;
import mem_ss_env_pkg::*;
import mem_ss_reg_pkg::*;
import mem_ss_seq_lib_pkg::*;

`include "mem_ss_test.svh"

endpackage: mem_ss_test_lib_pkg
