covergroup uart_cg_receive;

      option.per_instance = 1;

      selector: coverpoint trans.mode {


      bins addition0         = {'h080};
      bins subtraction0      = {'h081};
      bins multiplication0   = {'h082};
      bins division0         = {'h083};
      bins modulo_division0  = {'h084};
      bins logical_and0      = {'h085};
      bins logical_or0       = {'h086};
      bins logical_negation0 = {'h087};
      bins bitwise_negation0 = {'h088};
      bins bitwise_and0      = {'h089};
      bins bitwise_or0       = {'h08A};
      bins bitwise_xor0      = {'h08B};
      bins left_shift0       = {'h08C};
      bins right_shift0      = {'h08D};
      bins increment0        = {'h08E};
      bins decrement0        = {'h08F};
      bins add1tion0         = {'h090};
      bins subtract1on0      = {'h091};
      bins multiplicat1on0   = {'h092};
      bins divis1on0         = {'h093};
      bins modulo_divis1on0  = {'h094};
      bins log1cal_and0      = {'h095};
      bins log1cal_or0       = {'h096};
      bins log1cal_negation0 = {'h097};
      bins b1twise_negation0 = {'h098};
      bins b1twise_and0      = {'h099};
      bins b1twise_or0       = {'h09A};
      bins b1twise_xor0      = {'h09B};
      bins left_sh1ft0       = {'h09C};
      bins right_sh1ft0      = {'h09D};
      bins incremen10        = {'h09E};
      bins decremen10        = {'h09F};

      bins addition1         = {'h180};
      bins subtraction1      = {'h181};
      bins multiplication1   = {'h182};
      bins division1         = {'h183};
      bins modulo_division1  = {'h184};
      bins logical_and1      = {'h185};
      bins logical_or1       = {'h186};
      bins logical_negation1 = {'h187};
      bins bitwise_negation1 = {'h188};
      bins bitwise_and1      = {'h189};
      bins bitwise_or1       = {'h18A};
      bins bitwise_xor1      = {'h18B};
      bins left_shift1       = {'h18C};
      bins right_shift1      = {'h18D};
      bins increment1        = {'h18E};
      bins decrement1        = {'h18F};
      bins add1tion1         = {'h190};
      bins subtract1on1      = {'h191};
      bins multiplicat1on1   = {'h192};
      bins divis1on1         = {'h193};
      bins modulo_divis1on1  = {'h194};
      bins log1cal_and1      = {'h195};
      bins log1cal_or1       = {'h196};
      bins log1cal_negation1 = {'h197};
      bins b1twise_negation1 = {'h198};
      bins b1twise_and1      = {'h199};
      bins b1twise_or1       = {'h19A};
      bins b1twise_xor1      = {'h19B};
      bins left_sh1ft1       = {'h19C};
      bins right_sh1ft1      = {'h19D};
      bins incremen11        = {'h19E};
      bins decremen11        = {'h19F};

      bins addition2         = {'h280};
      bins subtraction2      = {'h281};
      bins multiplication2   = {'h282};
      bins division2         = {'h283};
      bins modulo_division2  = {'h284};
      bins logical_and2      = {'h285};
      bins logical_or2       = {'h286};
      bins logical_negation2 = {'h287};
      bins bitwise_negation2 = {'h288};
      bins bitwise_and2      = {'h289};
      bins bitwise_or2       = {'h28A};
      bins bitwise_xor2      = {'h28B};
      bins left_shift2       = {'h28C};
      bins right_shift2      = {'h28D};
      bins increment2        = {'h28E};
      bins decrement2        = {'h28F};
      bins add1tion2         = {'h290};
      bins subtract1on2      = {'h291};
      bins multiplicat1on2   = {'h292};
      bins divis1on2         = {'h293};
      bins modulo_divis1on2  = {'h294};
      bins log1cal_and2      = {'h295};
      bins log1cal_or2       = {'h296};
      bins log1cal_negation2 = {'h297};
      bins b1twise_negation2 = {'h298};
      bins b1twise_and2      = {'h299};
      bins b1twise_or2       = {'h29A};
      bins b1twise_xor2      = {'h29B};
      bins left_sh1ft2       = {'h29C};
      bins right_sh1ft2      = {'h29D};
      bins incremen12        = {'h29E};
      bins decremen12        = {'h29F};

      bins addition3         = {'h380};
      bins subtraction3      = {'h381};
      bins multiplication3   = {'h382};
      bins division3         = {'h383};
      bins modulo_division3  = {'h384};
      bins logical_and3      = {'h385};
      bins logical_or3       = {'h386};
      bins logical_negation3 = {'h387};
      bins bitwise_negation3 = {'h388};
      bins bitwise_and3      = {'h389};
      bins bitwise_or3       = {'h38A};
      bins bitwise_xor3      = {'h38B};
      bins left_shift3       = {'h38C};
      bins right_shift3      = {'h38D};
      bins increment3        = {'h38E};
      bins decrement3        = {'h38F};
      bins add1tion3         = {'h390};
      bins subtract1on3      = {'h391};
      bins multiplicat1on3   = {'h392};
      bins divis1on3         = {'h393};
      bins modulo_divis1on3  = {'h394};
      bins log1cal_and3      = {'h395};
      bins log1cal_or3       = {'h396};
      bins log1cal_negation3 = {'h397};
      bins b1twise_negation3 = {'h398};
      bins b1twise_and3      = {'h399};
      bins b1twise_or3       = {'h39A};
      bins b1twise_xor3      = {'h39B};
      bins left_sh1ft3       = {'h39C};
      bins right_sh1ft3      = {'h39D};
      bins incremen13        = {'h39E};
      bins decremen13        = {'h39F};


      option.at_least = 1;


    }   
 
endgroup 

