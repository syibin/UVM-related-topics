

wire            UART_SRX;   // UART serial input signal
wire            UART_STX;   // UART serial output signal
wire            UART_RTS;   // UART MODEM Request To Send
wire            UART_CTS;   // UART MODEM Clear To Send
wire            UART_DTR;   // UART MODEM Data Terminal Ready
wire            UART_DSR;   // UART MODEM Data Set Ready
wire            UART_RI;    // UART MODEM Ring Indicator
wire            UART_DCD;   // UART MODEM Data Carrier Detect

//UART internal
wire            UART_BAUD;  // UART baudrate output
wire            UART_INT;   // UART interrupt