package biquad_vseq_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

import apb_agent_pkg::*;
import signal_agent_pkg::*;
import biquad_reg_pkg::*;
import biquad_env_pkg::*;

`include "setup_coefficients.svh"
`include "biquad_vseq.svh"
`include "biquad_smoke_vseq.svh"

endpackage: biquad_vseq_pkg