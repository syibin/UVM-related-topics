covergroup uart_cg_loopback;
      option.per_instance = 1;
      selector: coverpoint trans.mode {

      bins addition0         = {'h0A0};
      bins subtraction0      = {'h0A1};
      bins multiplication0   = {'h0A2};
      bins division0         = {'h0A3};
      bins modulo_division0  = {'h0A4};
      bins logical_and0      = {'h0A5};
      bins logical_or0       = {'h0A6};
      bins logical_negation0 = {'h0A7};
      bins bitwise_negation0 = {'h0A8};
      bins bitwise_and0      = {'h0A9};
      bins bitwise_or0       = {'h0AA};
      bins bitwise_xor0      = {'h0AB};
      bins left_shift0       = {'h0AC};
      bins right_shift0      = {'h0AD};
      bins increment0        = {'h0AE};
      bins decrement0        = {'h0AF};
      bins add1tion0         = {'h0B0};
      bins subtract1on0      = {'h0B1};
      bins multiplicat1on0   = {'h0B2};
      bins divis1on0         = {'h0B3};
      bins modulo_divis1on0  = {'h0B4};
      bins log1cal_and0      = {'h0B5};
      bins log1cal_or0       = {'h0B6};
      bins log1cal_negation0 = {'h0B7};
      bins b1twise_negation0 = {'h0B8};
      bins b1twise_and0      = {'h0B9};
      bins b1twise_or0       = {'h0BA};
      bins b1twise_xor0      = {'h0BB};
      bins left_sh1ft0       = {'h0BC};
      bins right_sh1ft0      = {'h0BD};
      bins incremen10        = {'h0BE};
      bins decremen10        = {'h0BF};

      bins addition11        = {'h1A0};
      bins subtraction1      = {'h1A1};
      bins multiplication1   = {'h1A2};
      bins division1         = {'h1A3};
      bins modulo_division1  = {'h1A4};
      bins logical_and1      = {'h1A5};
      bins logical_or1       = {'h1A6};
      bins logical_negation1 = {'h1A7};
      bins bitwise_negation1 = {'h1A8};
      bins bitwise_and1      = {'h1A9};
      bins bitwise_or1       = {'h1AA};
      bins bitwise_xor1      = {'h1AB};
      bins left_shift1       = {'h1AC};
      bins right_shift1      = {'h1AD};
      bins increment1        = {'h1AE};
      bins decrement1        = {'h1AF};
      bins add1tion1         = {'h1B0};
      bins subtract1on1      = {'h1B1};
      bins multiplicat1on1   = {'h1B2};
      bins divis1on1         = {'h1B3};
      bins modulo_divis1on1  = {'h1B4};
      bins log1cal_and1      = {'h1B5};
      bins log1cal_or1       = {'h1B6};
      bins log1cal_negation1 = {'h1B7};
      bins b1twise_negation1 = {'h1B8};
      bins b1twise_and1      = {'h1B9};
      bins b1twise_or1       = {'h1BA};
      bins b1twise_xor1      = {'h1BB};
      bins left_sh1ft1       = {'h1BC};
      bins right_sh1ft1      = {'h1BD};
      bins incremen11        = {'h1BE};
      bins decremen11        = {'h1BF};
      
      bins addition2         = {'h2A0};
      bins subtraction2      = {'h2A1};
      bins multiplication2   = {'h2A2};
      bins division2         = {'h2A3};
      bins modulo_division2  = {'h2A4};
      bins logical_and2      = {'h2A5};
      bins logical_or2       = {'h2A6};
      bins logical_negation2 = {'h2A7};
      bins bitwise_negation2 = {'h2A8};
      bins bitwise_and2      = {'h2A9};
      bins bitwise_or2       = {'h2AA};
      bins bitwise_xor2      = {'h2AB};
      bins left_shift2       = {'h2AC};
      bins right_shift2      = {'h2AD};
      bins increment2        = {'h2AE};
      bins decrement2        = {'h2AF};
      bins add1tion2         = {'h2B0};
      bins subtract1on2      = {'h2B1};
      bins multiplicat1on2   = {'h2B2};
      bins divis1on2         = {'h2B3};
      bins modulo_divis1on2  = {'h2B4};
      bins log1cal_and2      = {'h2B5};
      bins log1cal_or2       = {'h2B6};
      bins log1cal_negation2 = {'h2B7};
      bins b1twise_negation2 = {'h2B8};
      bins b1twise_and2      = {'h2B9};
      bins b1twise_or2       = {'h2BA};
      bins b1twise_xor2      = {'h2BB};
      bins left_sh1ft2       = {'h2BC};
      bins right_sh1ft2      = {'h2BD};
      bins incremen12        = {'h2BE};
      bins decremen12        = {'h2BF};

      bins addition3         = {'h3A0};
      bins subtraction3      = {'h3A1};
      bins multiplication3   = {'h3A2};
      bins division3         = {'h3A3};
      bins modulo_division3  = {'h3A4};
      bins logical_and3      = {'h3A5};
      bins logical_or3       = {'h3A6};
      bins logical_negation3 = {'h3A7};
      bins bitwise_negation3 = {'h3A8};
      bins bitwise_and3      = {'h3A9};
      bins bitwise_or3       = {'h3AA};
      bins bitwise_xor3      = {'h3AB};
      bins left_shift3       = {'h3AC};
      bins right_shift3      = {'h3AD};
      bins increment3        = {'h3AE};
      bins decrement3        = {'h3AF};
      bins add1tion3         = {'h3B0};
      bins subtract1on3      = {'h3B1};
      bins multiplicat1on3   = {'h3B2};
      bins divis1on3         = {'h3B3};
      bins modulo_divis1on3  = {'h3B4};
      bins log1cal_and3      = {'h3B5};
      bins log1cal_or3       = {'h3B6};
      bins log1cal_negation3 = {'h3B7};
      bins b1twise_negation3 = {'h3B8};
      bins b1twise_and3      = {'h3B9};
      bins b1twise_or3       = {'h3BA};
      bins b1twise_xor3      = {'h3BB};
      bins left_sh1ft3       = {'h3BC};
      bins right_sh1ft3      = {'h3BD};
      bins incremen13        = {'h3BE};
      bins decremen13        = {'h3BF};

      option.at_least = 1;
    }    
endgroup 

