//
//------------------------------------------------------------------------------
//   Copyright 2010-2018 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------------------------

package dsp_con_pkg;

import uvm_pkg::*;
import interrupt_pkg::*;
`include "uvm_macros.svh"

`include "dsp_con_config.svh"
`include "dsp_con_seq_item.svh"
`include "dsp_con_sequencer.svh"
`include "dsp_con_driver.svh"
`include "dsp_con_agent.svh"
`include "dsp_con_seq.svh"
`include "dsp_con_test.svh"


endpackage: dsp_con_pkg
