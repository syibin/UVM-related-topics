//------------------------------------------------------------
//   Copyright 2010-2018 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------

package gpio_test_sequence_lib_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

import gpio_agent_pkg::*;
import gpio_env_pkg::*;
import gpio_bus_sequence_lib_pkg::*;

// This base class contains a body method implementation that assigns the
// sequencer handles to the actual sequences:
class gpio_virtual_sequence_base extends uvm_sequence #(uvm_sequence_item);

  `uvm_object_utils(gpio_virtual_sequence_base)

  function new(string name = "gpio_virtual_sequence_base");
    super.new(name);
  endfunction

  // env config object - needed to get to the wait_for_interrupt function
  gpio_env_config m_cfg;

  // Local handles for the sequencers
  gpio_sequencer gpi;
  gpio_sequencer aux;

  task body;
    // Check the sequencers
    if(gpi == null) begin
      `uvm_fatal("GPIO_SEQUENCERS", "The gpi sequencer handle is null - this simulation will fail");
    end

    // Getting access to the interrupt line
    if (m_cfg == null) begin
      `uvm_fatal("CONFIG_LOAD", "Configuration is null - this simulation will fail")
    end
  endtask: body

endclass: gpio_virtual_sequence_base

// Register test - checks reset and then R/W path
class reg_test_vseq extends gpio_virtual_sequence_base;

  `uvm_object_utils(reg_test_vseq)

  function new(string name = "reg_test_vseq");
    super.new(name);
  endfunction

  task body;
    //  check_reset_seq do_reset = check_reset_seq::type_id::create("do_reset");
    gpio_reg_rand reg_check = gpio_reg_rand::type_id::create("reg_check");
    gpio_seq init_gpio = gpio_seq::type_id::create("init_gpio");

    reg_check.m_cfg = m_cfg;

    // Get the virtual sequencer handles assigned
    super.body();

    // Initialise the GPI and AUX inputs to 0
    init_gpio.data = 0;
    if(aux != null) begin
      init_gpio.start(aux);
    end
    init_gpio.start(gpi);
    // Check the reset conditions
    //  do_reset.start(m_sequencer);
    reg_check.iterations = 200;
    reg_check.start(m_sequencer);
  endtask: body

endclass: reg_test_vseq

// GPIO Output path test
class GPO_test_vseq extends gpio_virtual_sequence_base;

  `uvm_object_utils(GPO_test_vseq)

  function new(string name = "GPO_test_vseq");
    super.new(name);
  endfunction

  task body();
    output_test_seq GP_OPs;
    gpio_rand_seq AUX_IPs;
    diag_outputs diag;
    aux_reg_seq AUX_reg;
    
    GP_OPs = output_test_seq::type_id::create("GP_OPs");
    AUX_IPs = gpio_rand_seq::type_id::create("AUX_IPs");
    diag = diag_outputs::type_id::create("diag");
    AUX_reg = aux_reg_seq::type_id::create("AUX_reg");

    GP_OPs.m_cfg = m_cfg;
    diag.m_cfg = m_cfg;
    AUX_reg.m_cfg = m_cfg;

    // Get the virtual sequencer handles assigned
    super.body();

    begin
      diag.start(m_sequencer);
      repeat(200) begin
        fork
          GP_OPs.start(m_sequencer);
          AUX_reg.start(m_sequencer);
        join
      end
    end

  endtask: body

endclass: GPO_test_vseq

// GPIO Input path test - including interrupts
class GPI_test_vseq extends gpio_virtual_sequence_base;

  `uvm_object_utils(GPI_test_vseq)

  function new(string name = "GPI_test_vseq");
    super.new(name);
  endfunction

  task body;
    gpio_isr ISR = gpio_isr::type_id::create("ISR");
    gpio_input_test_seq gpi_input_regs = gpio_input_test_seq::type_id::create("gpi_input_regs");
    gpio_rand_seq gpi_inputs = gpio_rand_seq::type_id::create("gpio_rand_seq");

    ISR.m_cfg = m_cfg;
    gpi_input_regs.m_cfg = m_cfg;

    super.body();

    fork
      gpi_inputs.start(gpi); // Forever
      begin // Setting up the GPI associated registers
        gpi_input_regs.iterations = 20000; // Repeat 100 times (Not enough)
        gpi_input_regs.start(m_sequencer);
      end
      begin // ISR
        forever begin
          m_cfg.wait_for_interrupt;
          ISR.start(m_sequencer);
        end
      end
    join_any

  endtask: body

endclass: GPI_test_vseq

endpackage: gpio_test_sequence_lib_pkg
