`define delay = 5
