//------------------------------------------------------------
//   Copyright 2010-2018 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------

module hdl_top;
  // pragma attribute hdl_top partition_module_xrtl

// PCLK and PRESETn
//
logic PCLK;
logic PRESETn;

wire[31:0] PADDR;
wire[31:0] PRDATA;
wire[31:0] PWDATA;
wire PWRITE;
wire PENABLE;
wire[31:0] PSEL;
wire PREADY;
wire PSLVERR;

//
// Instantiate the BFM interfaces:
//
apb_slave_driver_bfm  APB_slv_drv_bfm(.PCLK(PCLK),
                                      .PRESETn(PRESETn),
                                      .PADDR(PADDR),
                                      .PRDATA(PRDATA),
                                      .PWDATA(PWDATA),
                                      .PSEL(PSEL),
                                      .PENABLE(PENABLE),
                                      .PWRITE(PWRITE),
                                      .PREADY(PREADY),
                                      .PSLVERR(PSLVERR));
                                      
apb_slave_monitor_bfm APB_slv_mon_bfm(.PCLK(PCLK),
                                      .PRESETn(PRESETn),
                                      .PADDR(PADDR),
                                      .PRDATA(PRDATA),
                                      .PWDATA(PWDATA),
                                      .PSEL(PSEL),
                                      .PENABLE(PENABLE),
                                      .PWRITE(PWRITE),
                                      .PREADY(PREADY),
                                      .PSLVERR(PSLVERR));

    
apb3_wlm_host master (.pclk(PCLK), 
                      .presetn(PRESETn), 
                      .paddr(PADDR), 
                      .psel(PSEL[0]), 
                      .penable(PENABLE),
                      .pwrite(PWRITE), 
                      .pwdata(PWDATA), 
                      .prdata(PRDATA), 
                      .pready(PREADY), 
                      .pslverr(PSLVERR));


// UVM initial block:
// Virtual interface wrapping 
initial begin //tbx vif_binding_block
  import uvm_pkg::uvm_config_db;
  uvm_config_db #(virtual apb_slave_driver_bfm) ::set(null, "uvm_test_top", "APB_slv_drv_bfm", APB_slv_drv_bfm);
  uvm_config_db #(virtual apb_slave_monitor_bfm) ::set(null, "uvm_test_top", "APB_slv_mon_bfm", APB_slv_mon_bfm);
end

assign PSEL[15:1] = 'b1;
//
// Clock and reset initial block:
//
initial begin
  PCLK = 0;
  PRESETn = 0;
  repeat(8) begin
    #10ns PCLK = ~PCLK;
  end
  PRESETn = 1;
  forever begin
    #10ns PCLK = ~PCLK;
  end
end

endmodule: hdl_top
