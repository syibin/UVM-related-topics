wait(uif.interrupt[2]);
if(uif.interrupt[2] & ins_errors[0]) begin : FERR

    wait(uif.interrupt[2]);
    $display("\033[1;31mError Interrupt Has Been Asserted. Time : %t\033[0m", $realtime);

    do  begin
        reg_access( `UART_BASE_ADDRESS + `UART_STATUS_REGISTER,
                    REG_RD,
                    32'h0,
                    4'h0,
                    read_data,
                    error
                  );
        end
    while(!read_data[2]);

    if(!read_data[2]) begin

      $display("\033[1;31mFraming error was not detected during RECEIVE_FRAMING_ERROR test\033[0m");
      print_test_result("FAILED");
      $finish(2);

    end

    if(!symbol[8]) begin

      $display("\033[1;31mIllegaly detected framing error during data receiption @%t. Testbench didn't generate this error\033[0m", $time);
      print_test_result("FAILED");
      $finish(2);

    end

    else if(symbol[8]) begin
      $display("\033[1;32mDetected framing error correctly generated by testbench @%t\033[0m", $time);

      reg_access( `UART_BASE_ADDRESS + `UART_RXBUF_REGISTER,
                  REG_RD,
                  32'h0,
                  4'h0,
                  read_data,
                  error
                );
    end

end : FERR

else begin : FERR_N

      $display("\033[1;31mWRONG!!Error Interrupt hasn't been Asserted!! FERR @Time %t\033[0m", $realtime);
      //$finish;

end : FERR_N