package spi_agent_pkg;
  
  import uvm_pkg::*;
    
  `include "uvm_macros.svh"
  
  `include "C:\\Users\\Boolman\\Desktop\\ankasys_project\\agent\\spi_item.svh"
  `include "C:\\Users\\Boolman\\Desktop\\ankasys_project\\agent\\spi_test_config.svh"
  `include "C:\\Users\\Boolman\\Desktop\\ankasys_project\\agent\\spi_sequence.svh"
  `include "C:\\Users\\Boolman\\Desktop\\ankasys_project\\agent\\spi_sequencer.svh"
  `include "C:\\Users\\Boolman\\Desktop\\ankasys_project\\agent\\spi_monitor.svh"
  `include "C:\\Users\\Boolman\\Desktop\\ankasys_project\\agent\\spi_driver.svh"
  `include "C:\\Users\\Boolman\\Desktop\\ankasys_project\\agent\\spi_agent.svh"

endpackage