//------------------------------------------------------------
//   Copyright 2010-2018 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------

module hdl_top;

`include "gpio_defines.v"
`include "timescale.v"

// PCLK and PRESETn
//
logic PCLK;
logic PRESETn;

//
// Instantiate the pin interfaces:
//
apb_if APB(PCLK, PRESETn);   // APB interface
gpio_if GPO();  // GPO Output
gpio_if GPOE(); // GPO Output Enable
gpio_if GPI();  // GPI Input
gpio_if AUX();  // GPO Auxillary Input
intr_if INTR();   // Interrupt

//
// Instantiate the BFM interfaces:
//
apb_monitor_bfm APB_mon_bfm(
   .PCLK    (APB.PCLK),
   .PRESETn (APB.PRESETn),
   .PADDR   (APB.PADDR),
   .PRDATA  (APB.PRDATA),
   .PWDATA  (APB.PWDATA),
   .PSEL    (APB.PSEL),
   .PENABLE (APB.PENABLE),
   .PWRITE  (APB.PWRITE),
   .PREADY  (APB.PREADY)
);
apb_driver_bfm  APB_drv_bfm(
   .PCLK    (APB.PCLK),
   .PRESETn (APB.PRESETn),
   .PADDR   (APB.PADDR),
   .PRDATA  (APB.PRDATA),
   .PWDATA  (APB.PWDATA),
   .PSEL    (APB.PSEL),
   .PENABLE (APB.PENABLE),
   .PWRITE  (APB.PWRITE),
   .PREADY  (APB.PREADY)
);
gpio_monitor_bfm GPO_mon_bfm(
   .clk     (GPO.clk),
   .gpio    (GPO.gpio),
   .ext_clk (GPO.ext_clk)
);
//gpio_driver_bfm  GPO_drv_bfm(
//   .clk     (GPO.clk),
//   .gpio    (GPO.gpio),
//   .ext_clk (GPO.ext_clk)
//);
gpio_monitor_bfm GPOE_mon_bfm(
   .clk     (GPOE.clk),
   .gpio    (GPOE.gpio),
   .ext_clk (GPOE.ext_clk)
);
//gpio_driver_bfm  GPOE_drv_bfm(
//   .clk     (GPOE.clk),
//   .gpio    (GPOE.gpio),
//   .ext_clk (GPOE.ext_clk)
//);
gpio_monitor_bfm GPI_mon_bfm(
   .clk     (GPI.clk),
   .gpio    (GPI.gpio),
   .ext_clk (GPI.ext_clk)
);
gpio_driver_bfm  GPI_drv_bfm(
   .clk     (GPI.clk),
   .gpio    (GPI.gpio),
   .ext_clk (GPI.ext_clk)
);
gpio_monitor_bfm AUX_mon_bfm(
   .clk     (AUX.clk),
   .gpio    (AUX.gpio),
   .ext_clk (AUX.ext_clk)
);
gpio_driver_bfm  AUX_drv_bfm(
   .clk     (AUX.clk),
   .gpio    (AUX.gpio),
   .ext_clk (AUX.ext_clk)
);


// DUT
gpio_top DUT(
  // APB Interface:
  .PCLK(PCLK),
  .PRESETN(PRESETn),
  .PSEL(APB.PSEL[0]),
  .PADDR(APB.PADDR[7:0]),
  .PWDATA(APB.PWDATA),
  .PRDATA(APB.PRDATA),
  .PENABLE(APB.PENABLE),
  .PREADY(APB.PREADY),
  .PSLVERR(),
  .PWRITE(APB.PWRITE),
  // Interrupt output
  .IRQ(INTR.IRQ),
`ifdef GPIO_AUX_IMPLEMENT
  // Auxiliary inputs interface
  .aux_i(AUX.gpio),
`endif //  GPIO_AUX_IMPLEMENT
  // External GPIO Interface
  .ext_pad_i(GPI.gpio),
  .ext_pad_o(GPO.gpio),
  .ext_padoe_o(GPOE.gpio)
`ifdef GPIO_CLKPAD
  , .clk_pad_i(GPI.ext_clk)
`endif
);

// UVM initial block:
// Virtual interface wrapping & run_test()
initial begin //tbx vif_binding_block
  import uvm_pkg::uvm_config_db;
  uvm_config_db #(virtual apb_monitor_bfm)::set(null, "uvm_test_top", "APB_mon_bfm", APB_mon_bfm);
  uvm_config_db #(virtual apb_driver_bfm) ::set(null, "uvm_test_top", "APB_drv_bfm", APB_drv_bfm);
  uvm_config_db #(virtual gpio_monitor_bfm)::set(null, "uvm_test_top", "GPO_mon_bfm", GPO_mon_bfm);
//  uvm_config_db #(virtual gpio_driver_bfm) ::set(null, "uvm_test_top", "GPO_drv_bfm", GPO_drv_bfm);
  uvm_config_db #(virtual gpio_monitor_bfm)::set(null, "uvm_test_top", "GPOE_mon_bfm", GPOE_mon_bfm);
//  uvm_config_db #(virtual gpio_driver_bfm) ::set(null, "uvm_test_top", "GPOE_drv_bfm", GPOE_drv_bfm);
  uvm_config_db #(virtual gpio_monitor_bfm)::set(null, "uvm_test_top", "GPI_mon_bfm", GPI_mon_bfm);
  uvm_config_db #(virtual gpio_driver_bfm) ::set(null, "uvm_test_top", "GPI_drv_bfm", GPI_drv_bfm);
  uvm_config_db #(virtual gpio_monitor_bfm)::set(null, "uvm_test_top", "AUX_mon_bfm", AUX_mon_bfm);
  uvm_config_db #(virtual gpio_driver_bfm) ::set(null, "uvm_test_top", "AUX_drv_bfm", AUX_drv_bfm);
  uvm_config_db #(virtual intr_if)::set(null, "uvm_test_top", "INTR_vif", INTR);
end

//
// Clock and reset initial block:
//
initial begin
  PCLK = 0;
  forever #10ns PCLK = ~PCLK;
end
initial begin 
  PRESETn = 0;
  repeat(4) @(posedge PCLK);
  PRESETn = 1;
end

// Clock assignments:
assign GPO.clk = PCLK;
assign GPOE.clk = PCLK;
assign AUX.clk = PCLK;
assign GPI.clk = PCLK;

endmodule: hdl_top
