//------------------------------------------------------------
//   Copyright 2010-2018 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//   
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//   
//       http://www.apache.org/licenses/LICENSE-2.0
//   
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------

// hvl_top level module for rtl alu
module hvl_top();
import uvm_pkg::*;
import alu_tb_pkg::*;

 initial begin
     // start with default "test" (using std_stim_group) 
     // override this with plusarg UVM_TESTNAME
  run_test("test_std_stim_gen");
 end
  
endmodule : hvl_top
