//*****************************************************************************
// This test checks data receiption with ability of errors insertion by
// testbench
//
// The sequence of steps is:
//
// 1) Wait for the end of reset, then wait 10 clocks
// 2) Program MODE and INTC Registers
// 3) Testbench in a loop generates activity on rxd line of DUT to send a
//    character
// 4) Testbench waits for interrupt and handle it according to the test
//    configuration (existense of errors insertion)
//*****************************************************************************

print_test_config( `UART_STATUS_REGISTER,
                   mode,
                   interrupts_config,
                   `CHARACTER_NUM
                 );


wait(rst_n);
repeat(10) @(posedge clk);


//program MODE register
reg_access( `UART_BASE_ADDRESS + `UART_MODE_REGISTER,
            REG_WR,
            mode,
            4'h3,
            read_data,
            error
          );

if(error) begin
  $display("Error occured during setting up UART's operation mode, address is 32'h%h, data is 32'h%h, byte enable is",
           `UART_BASE_ADDRESS + 32'h8, mode, 4'h1
          );
  $finish(2);
end

//program INTC Register
reg_access( `UART_BASE_ADDRESS + `UART_INTC_REGISTER,
            REG_WR,
            {29'b0, interrupts_config},
            4'h1,
            read_data,
            error
          );


//repeat CHARACTER_NUM symbols receiption
if(!mode[9]) repeat (`CHARACTER_NUM) begin : uart_rx_single_bytes

  send_error = $urandom_range(8,0);
  $display("send_error = %0h", send_error);


  if(|send_error) send_uart_char( ins_errors[1],
                                  ins_errors[0],
                                  mode
                                );
   else           send_uart_char( 1'b0,
                                  1'b0,
                                  mode
                                );

  wait(interrupt);

  reg_access( `UART_BASE_ADDRESS + `UART_INTF_REGISTER,
              REG_RD,
              32'h0,
              4'h0,
              read_data,
              error
            );

  intf = read_data;


  reg_access( `UART_BASE_ADDRESS + `UART_STATUS_REGISTER,
              REG_RD,
              32'h0,
              4'h0,
              read_data,
              error
            );

  if(intf[2] & ins_errors[1] & (|send_error)) begin


    if(!read_data[3]) begin
      $display("Parity error was not detected during RECEIVE_PARITY_ERROR test");
      print_test_result("FAILED");
      $finish(2);
    end

    symbol = rx_data_queue.pop_front();
    if(!symbol[9]) begin
      $display("Illegaly detected parity error during data receiption @%t. Testbench didn't generate this error", $time);
      print_test_result("FAILED");
      $finish(2);
    end
    else begin
      $display("Detected parity error correctly generated by testbench @%t", $time);

      if(!read_data[2]) begin
        reg_access( `UART_BASE_ADDRESS + `UART_RXBUF_REGISTER,
                    REG_RD,
                    32'h0,
                    4'h0,
                    read_data,
                    error
                  );
      end

    end

  end


  if(intf[2] & ins_errors[0] & (|send_error)) begin


    reg_access( `UART_BASE_ADDRESS + `UART_STATUS_REGISTER,
                REG_RD,
                32'h0,
                4'h0,
                read_data,
                error
              );


    if(!read_data[2]) begin
      $display("Framing error was not detected during RECEIVE_FRAMING_ERROR test");
      print_test_result("FAILED");
      $finish(2);
    end

    if(!read_data[3]) symbol = rx_data_queue.pop_front();
    if(!symbol[8]) begin
      $display("Illegaly detected framing error during data receiption @%t. Testbench didn't generate this error", $time);
      print_test_result("FAILED");
      $finish(2);
    end
    else begin
      $display("Detected framing error correctly generated by testbench @%t", $time);

      reg_access( `UART_BASE_ADDRESS + `UART_RXBUF_REGISTER,
                  REG_RD,
                  32'h0,
                  4'h0,
                  read_data,
                  error
                );
    end

  end


  if(intf[0]) begin
    $display("Illegal interrupt set");
    print_test_result("FAILED");
    $finish(2);
  end

  symbol = rx_data_queue.pop_front();


  if(intf[1] & (!(|ins_errors) | !(|send_error))) begin : handle_rx_int

    //read data from RXBUF
    reg_access( `UART_BASE_ADDRESS + `UART_RXBUF_REGISTER,
                REG_RD,
                32'h0,
                4'h0,
                read_data,
                error
              );

    //check if received data is correct (the same as it was sent)
    if(symbol[7:0] != read_data[7:0]) begin
      $display("Received character doesn't match the character sent by testbench! Received \"%s\", sent \"%s\"", read_data[7:0], symbol);
      print_test_result("FAILED");
      $finish(2);
    end
    else $display("Received character matches the character sent by testbench. Received \"%s\", sent \"%s\"", read_data[7:0], symbol);

  end : handle_rx_int

  if(intf[1] & !intf[2] & (|ins_errors)) begin

    //read data from RXBUF
    reg_access( `UART_BASE_ADDRESS + `UART_RXBUF_REGISTER,
                REG_RD,
                32'h0,
                4'h0,
                read_data,
                error
              );
  end


  //clean interrupt flags
  reg_access( `UART_BASE_ADDRESS + `UART_INTF_REGISTER,
              REG_WR,
              {29'b0, 3'b111},
              4'h1,
              read_data,
              error
            );



end : uart_rx_single_bytes

else if(mode[9:8] == 2'b10) begin : uart_rx_triple_byte

  if((`CHARACTER_NUM / 3 == 0) | (`CHARACTER_NUM % 3 != 0)) begin
    $display("Test scenario is not valid. Controller programmed to generate interrupt after reception of 3 bytes, but CHARACTER_NUM parameter is not an integer number of 3-byte portions");
    $finish(2);
  end

  else repeat(`CHARACTER_NUM / 3) begin : rcv_3b_chunk

    //send 3 characters to UART Receiver
    repeat(3) begin

      if(|send_error) send_uart_char( ins_errors[1],
                                      ins_errors[0],
                                      mode
                                    );
      else            send_uart_char( 1'b0,
                                      1'b0,
                                      mode
                                    );

      repeat(5) @(posedge clk);

    end

    wait(interrupt);

    reg_access( `UART_BASE_ADDRESS + `UART_INTF_REGISTER,
                REG_RD,
                32'h0,
                4'h0,
                read_data,
                error
              );

    intf = read_data;


    reg_access( `UART_BASE_ADDRESS + `UART_STATUS_REGISTER,
                REG_RD,
                32'h0,
                4'h0,
                read_data,
                error
              );

    symbol = rx_data_queue.pop_front();


    if(intf[1] & (!(|ins_errors) | !(|send_error))) begin : handle_rx3b_int

      //read data from RXBUF
      reg_access( `UART_BASE_ADDRESS + `UART_RXBUF_REGISTER,
                  REG_RD,
                  32'h0,
                  4'h0,
                  read_data,
                  error
                );

      //check if received data is correct (the same as it was sent)
      if(symbol[23:0] != read_data[23:0]) begin
        $display("Received character doesn't match the character sent by testbench! Received \"%s\", sent \"%s\"", read_data[23:0], symbol);
        print_test_result("FAILED");
        $finish(2);
      end
      else $display("Received character matches the character sent by testbench. Received \"%s\", sent \"%s\"", read_data[23:0], symbol);

    end : handle_rx3b_int

  end : rcv_3b_chunk


  //clean interrupt flags
  reg_access( `UART_BASE_ADDRESS + `UART_INTF_REGISTER,
              REG_WR,
              {29'b0, 3'b111},
              4'h1,
              read_data,
              error
            );


end : uart_rx_triple_byte


print_test_result("PASSED");
$finish(2);


