package spi_test_pkg;
  
  import uvm_pkg::*;
  import spi_agent_pkg::*;
    
  `include "uvm_macros.svh"
  
  `include "C:\\Users\\Boolman\\Desktop\\ankasys_project\\spi_env.svh"
  `include "C:\\Users\\Boolman\\Desktop\\ankasys_project\\spi_test.svh"


endpackage