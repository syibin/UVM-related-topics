`ifdef r128a32_25um
`else
`define r128a32_25um
`include "ram128x18_25um.v"
/************************************************************************
** File : r128a32_25um.v
** Design Date: June 9, 1998
** Creation Date: Mon Apr 15 15:16:35 2002

** Created By SpDE Version: SpDE 9.2 Release Build8
** Author: Robert Maul, QuickLogic Corporation,
** Copyright (C) 1998, Customers of QuickLogic may copy and modify this
** file for use in designing QuickLogic devices only.
** Description : This file is autogenerated RTL code that describes the
** connectivity of cascaded RAM blocks (RAM banks) using QuickLogic's
** RAM block resources.
************************************************************************/

module r128a32_25um(wa,ra,wd,rd,we,wclk);

// inputs: =wa[6:0]=,=ra[6:0]=,=wd[31:0]=,we,wclk
// outputs: =rd[31:0]=

input we;
input wclk;
input [6:0] wa;
input [6:0] ra;
input [31:0] wd;
output [31:0] rd;
supply0 GND;
supply1 VCC;
RAM128X18_25UM r128a32_25umI1 (.WA(wa),.RA(ra),.WD(wd[31:14]),.RD(rd[31:14]),
  .WE(we),.RE(GND),.WCLK(wclk),.RCLK(GND),.ASYNCRD(VCC));
RAM128X18_25UM r128a32_25umI2 (.WA(wa),.RA(ra),.WD({wd[13],wd[12],wd[11],wd[10],wd[9],wd[8],wd[7],wd[6],wd[5],wd[4],wd[3],wd[2],wd[1],wd[0], GND, GND, GND, GND}),.RD({rd[13],rd[12],rd[11],rd[10],rd[9],rd[8],rd[7],rd[6],rd[5],rd[4],rd[3],rd[2],rd[1],rd[0], dummy0, dummy1, dummy2, dummy3}),
  .WE(we),.RE(GND),.WCLK(wclk),.RCLK(GND),.ASYNCRD(VCC));
endmodule
`endif
