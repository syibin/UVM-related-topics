`include "./uart_xtn.sv"
`include "./uart_tx_sequencer.sv"
`include "./uart_tx_vsequencer.sv"
`include "./uart_tx_driver.sv"
`include "./uart_tx_monitor.sv"
`include "./uart_dut_monitor.sv"
`include "./uart_tx_agent.sv"
`include "./uart_dut_agent.sv"
`include "./uart_tx_uvc.sv"
`include "./../top/uart_tx_sb.sv"
`include "./../top/uart_tb.sv"
`include "./../sequences/uart_seqs.sv"
`include "./../sequences/uart_vseqs.sv"
