/* Verilog Model Created from SCS Schematic macros.sch */
/* From: 	Sandya@quicklogic.com */
/* Date:	August 31, 2001 */
/* Revision: 1.1 */
/* 8/31/01  Added Synthesis attributes (syn_isclock=1 and black_box_tri_pin)
for rev1.1 (sandya) */
/* If you are simulating a 0.25 micron device, you should copy 
'macros-25.v' to 'macros.v' before starting simulation. */
/* If you are simulating pre-0.25 micron devices, you should copy 
'macros-original.v' to 'macros.v' before starting simulation. */
/* Automatically generated by hvveri version 9.1 */

`timescale 1ns/1ns  
`define LOGIC   1 
`define BIDIR   2 
`define INCELL  3 
`define CLOCK   4 
`define HSCK    5 
`define CLOCKB  6 
`define ESPXCLKIN  7 
`define HSCKMUX 8 
`define IOCONTROL 9 



`ifdef upflct32
`else
`define upflct32
module upflct32( CLK , CLR, D, LOAD, Q );
input CLK  /* synthesis syn_isclock=1 */;
input CLR  /* synthesis syn_isclock=1 */;
 input [0:31] D;
input LOAD;
 output [0:31] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;

upflct4a QL11 ( .CLK(CLK), .CLR(CLR), .D({ D[0:3] }), .LOAD(LOAD), .Q({ Q[0:3] }),
             .RCO(N_14) );
upflct4b QL10 ( .CLK(CLK), .CLR(CLR), .D({ D[20:23] }), .ENP(N_7), .ENT(N_11),
             .LOAD(LOAD), .Q({ Q[20:23] }), .RCO(N_12) );
upflct4b QL9 ( .CLK(CLK), .CLR(CLR), .D({ D[24:27] }), .ENP(N_4), .ENT(N_12),
            .LOAD(LOAD), .Q({ Q[24:27] }), .RCO(N_13) );
upflct4b QL8 ( .CLK(CLK), .CLR(CLR), .D({ D[16:19] }), .ENP(N_3), .ENT(N_10),
            .LOAD(LOAD), .Q({ Q[16:19] }), .RCO(N_11) );
upflct4b QL7 ( .CLK(CLK), .CLR(CLR), .D({ D[12:15] }), .ENP(N_6), .ENT(N_9),
            .LOAD(LOAD), .Q({ Q[12:15] }), .RCO(N_10) );
upflct4b QL6 ( .CLK(CLK), .CLR(CLR), .D({ D[8:11] }), .ENP(N_2), .ENT(N_8),
            .LOAD(LOAD), .Q({ Q[8:11] }), .RCO(N_9) );
upflct4b QL5 ( .CLK(CLK), .CLR(CLR), .D({ D[4:7] }), .ENP(N_5), .ENT(N_14),
            .LOAD(LOAD), .Q({ Q[4:7] }), .RCO(N_8) );
upflct4c QL4 ( .CLK(CLK), .CLR(CLR), .D({ D[28:31] }), .ENP(N_1), .ENT(N_13),
            .LOAD(LOAD), .Q({ Q[28:31] }) );
upflcar2 QL3 ( .ACO1(N_6), .ACO2(N_3), .CLK(CLK), .CLR(CLR), .D({ D[0:1] }),
            .LOAD(LOAD) );
upflcar2 QL2 ( .ACO1(N_5), .ACO2(N_2), .CLK(CLK), .CLR(CLR), .D({ D[0:1] }),
            .LOAD(LOAD) );
upflcar3 QL1 ( .ACO1(N_7), .ACO2(N_4), .ACO3(N_1), .CLK(CLK), .CLR(CLR),
            .D({ D[0:1] }), .LOAD(LOAD) );

endmodule // upflct32

`endif

`ifdef upfxct8
`else
`define upfxct8
module upfxct8( CLK , CLR, D, EN, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:7] D;
input EN, LOAD;
 output [0:7] Q;
wire N_1;
wire N_2;

upfxcar1 QL3 ( .ACO1(N_1), .CLK(CLK), .CLR(CLR), .D({ D[0:1] }), .ENG(EN),
            .LOAD(LOAD), .Q({ Q[0:1] }) );
upfxct4c QL2 ( .CLK(CLK), .CLR(CLR), .D({ D[4:7] }), .ENG(EN), .ENP(N_1),
            .ENT(N_2), .LOAD(LOAD), .Q({ Q[4:7] }) );
upfxct4a QL1 ( .CLK(CLK), .CLR(CLR), .D({ D[0:3] }), .ENG(EN), .LOAD(LOAD),
            .Q({ Q[0:3] }), .RCO(N_2) );

endmodule // upfxct8

`endif

`ifdef upfxct4
`else
`define upfxct4
module upfxct4( CLK , CLR, D, EN, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:3] D;
input EN, LOAD;
 output [0:3] Q;
supply0 GND;

upfxct4c QL1 ( .CLK(CLK), .CLR(CLR), .D({ D[0:3] }), .ENG(EN), .ENP(GND),
            .ENT(GND), .LOAD(LOAD), .Q({ Q[0:3] }) );

endmodule // upfxct4

`endif

`ifdef upfxct32
`else
`define upfxct32
module upfxct32( CLK , CLR, D, EN, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:31] D;
input EN, LOAD;
 output [0:31] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;

upfxct4c QL11 ( .CLK(CLK), .CLR(CLR), .D({ D[28:31] }), .ENG(EN), .ENP(N_1),
             .ENT(N_4), .LOAD(LOAD), .Q({ Q[28:31] }) );
upfxcar3 QL10 ( .ACO1(N_11), .ACO2(N_10), .ACO3(N_9), .CLK(CLK), .CLR(CLR),
             .D({ D[0:1] }), .ENG(EN), .LOAD(LOAD), .Q({ Q[0:1] }) );
upfxcar2 QL9 ( .ACO1(N_2), .ACO2(N_1), .CLK(CLK), .CLR(CLR), .D({ D[0:1] }),
            .ENG(EN), .LOAD(LOAD) );
upfxcar2 QL8 ( .ACO1(N_6), .ACO2(N_5), .CLK(CLK), .CLR(CLR), .D({ D[0:1] }),
            .ENG(EN), .LOAD(LOAD) );
upfxct4a QL7 ( .CLK(CLK), .CLR(CLR), .D({ D[0:3] }), .ENG(EN), .LOAD(LOAD),
            .Q({ Q[0:3] }), .RCO(N_14) );
upfxct4b QL6 ( .CLK(CLK), .CLR(CLR), .D({ D[24:27] }), .ENG(EN), .ENP(N_2),
            .ENT(N_3), .LOAD(LOAD), .Q({ Q[24:27] }), .RCO(N_4) );
upfxct4b QL5 ( .CLK(CLK), .CLR(CLR), .D({ D[20:23] }), .ENG(EN), .ENP(N_5),
            .ENT(N_8), .LOAD(LOAD), .Q({ Q[20:23] }), .RCO(N_3) );
upfxct4b QL4 ( .CLK(CLK), .CLR(CLR), .D({ D[16:19] }), .ENG(EN), .ENP(N_6),
            .ENT(N_7), .LOAD(LOAD), .Q({ Q[16:19] }), .RCO(N_8) );
upfxct4b QL3 ( .CLK(CLK), .CLR(CLR), .D({ D[12:15] }), .ENG(EN), .ENP(N_9),
            .ENT(N_13), .LOAD(LOAD), .Q({ Q[12:15] }), .RCO(N_7) );
upfxct4b QL2 ( .CLK(CLK), .CLR(CLR), .D({ D[8:11] }), .ENG(EN), .ENP(N_10),
            .ENT(N_12), .LOAD(LOAD), .Q({ Q[8:11] }), .RCO(N_13) );
upfxct4b QL1 ( .CLK(CLK), .CLR(CLR), .D({ D[4:7] }), .ENG(EN), .ENP(N_11),
            .ENT(N_14), .LOAD(LOAD), .Q({ Q[4:7] }), .RCO(N_12) );

endmodule // upfxct32

`endif

`ifdef upfxct24
`else
`define upfxct24
module upfxct24( CLK , CLR, D, EN, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:23] D;
input EN, LOAD;
 output [0:23] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;

upfxct4c QL8 ( .CLK(CLK), .CLR(CLR), .D({ D[20:23] }), .ENG(EN), .ENP(N_1),
            .ENT(N_3), .LOAD(LOAD), .Q({ Q[20:23] }) );
upfxcar3 QL7 ( .ACO1(N_7), .ACO2(N_6), .ACO3(N_5), .CLK(CLK), .CLR(CLR),
            .D({ D[0:1] }), .ENG(EN), .LOAD(LOAD), .Q({ Q[0:1] }) );
upfxcar2 QL6 ( .ACO1(N_2), .ACO2(N_1), .CLK(CLK), .CLR(CLR), .D({ D[0:1] }),
            .ENG(EN), .LOAD(LOAD) );
upfxct4a QL5 ( .CLK(CLK), .CLR(CLR), .D({ D[0:3] }), .ENG(EN), .LOAD(LOAD),
            .Q({ Q[0:3] }), .RCO(N_10) );
upfxct4b QL4 ( .CLK(CLK), .CLR(CLR), .D({ D[16:19] }), .ENG(EN), .ENP(N_2),
            .ENT(N_4), .LOAD(LOAD), .Q({ Q[16:19] }), .RCO(N_3) );
upfxct4b QL3 ( .CLK(CLK), .CLR(CLR), .D({ D[12:15] }), .ENG(EN), .ENP(N_5),
            .ENT(N_9), .LOAD(LOAD), .Q({ Q[12:15] }), .RCO(N_4) );
upfxct4b QL2 ( .CLK(CLK), .CLR(CLR), .D({ D[8:11] }), .ENG(EN), .ENP(N_6),
            .ENT(N_8), .LOAD(LOAD), .Q({ Q[8:11] }), .RCO(N_9) );
upfxct4b QL1 ( .CLK(CLK), .CLR(CLR), .D({ D[4:7] }), .ENG(EN), .ENP(N_7),
            .ENT(N_10), .LOAD(LOAD), .Q({ Q[4:7] }), .RCO(N_8) );

endmodule // upfxct24

`endif

`ifdef upfxct16
`else
`define upfxct16
module upfxct16( CLK , CLR, D, EN, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:15] D;
input EN, LOAD;
 output [0:15] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;

upfxcar3 QL5 ( .ACO1(N_3), .ACO2(N_2), .ACO3(N_1), .CLK(CLK), .CLR(CLR),
            .D({ D[0:1] }), .ENG(EN), .LOAD(LOAD), .Q({ Q[0:1] }) );
upfxct4c QL4 ( .CLK(CLK), .CLR(CLR), .D({ D[12:15] }), .ENG(EN), .ENP(N_1),
            .ENT(N_5), .LOAD(LOAD), .Q({ Q[12:15] }) );
upfxct4b QL3 ( .CLK(CLK), .CLR(CLR), .D({ D[8:11] }), .ENG(EN), .ENP(N_2),
            .ENT(N_4), .LOAD(LOAD), .Q({ Q[8:11] }), .RCO(N_5) );
upfxct4b QL2 ( .CLK(CLK), .CLR(CLR), .D({ D[4:7] }), .ENG(EN), .ENP(N_3),
            .ENT(N_6), .LOAD(LOAD), .Q({ Q[4:7] }), .RCO(N_4) );
upfxct4a QL1 ( .CLK(CLK), .CLR(CLR), .D({ D[0:3] }), .ENG(EN), .LOAD(LOAD),
            .Q({ Q[0:3] }), .RCO(N_6) );

endmodule // upfxct16

`endif

`ifdef upflct8
`else
`define upflct8
module upflct8( CLK , CLR, D, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:7] D;
input LOAD;
 output [0:7] Q;
wire N_1;
supply0 GND;

upflcar1 QL3 ( .ACO1(N_1), .CLK(CLK), .CLR(CLR), .D({ D[0:3] }), .LOAD(LOAD),
            .Q({ Q[0:3] }) );
upflct4c QL2 ( .CLK(CLK), .CLR(CLR), .D({ D[0:3] }), .ENP(GND), .ENT(GND),
            .LOAD(LOAD), .Q({ Q[0:3] }) );
upflct4c QL1 ( .CLK(CLK), .CLR(CLR), .D({ D[4:7] }), .ENP(N_1), .ENT(GND),
            .LOAD(LOAD), .Q({ Q[4:7] }) );

endmodule // upflct8

`endif

`ifdef upflct4
`else
`define upflct4
module upflct4( CLK , CLR, D, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:3] D;
input LOAD;
 output [0:3] Q;
supply0 GND;

upflct4c QL1 ( .CLK(CLK), .CLR(CLR), .D({ D[0:3] }), .ENP(GND), .ENT(GND),
            .LOAD(LOAD), .Q({ Q[0:3] }) );

endmodule // upflct4

`endif

`ifdef upflct24
`else
`define upflct24
module upflct24( CLK , CLR, D, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:23] D;
input LOAD;
 output [0:23] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;

upflct4a QL8 ( .CLK(CLK), .CLR(CLR), .D({ D[0:3] }), .LOAD(LOAD), .Q({ Q[0:3] }),
            .RCO(N_10) );
upflct4b QL7 ( .CLK(CLK), .CLR(CLR), .D({ D[16:19] }), .ENP(N_2), .ENT(N_4),
            .LOAD(LOAD), .Q({ Q[16:19] }), .RCO(N_5) );
upflct4b QL6 ( .CLK(CLK), .CLR(CLR), .D({ D[12:15] }), .ENP(N_3), .ENT(N_9),
            .LOAD(LOAD), .Q({ Q[12:15] }), .RCO(N_4) );
upflct4b QL5 ( .CLK(CLK), .CLR(CLR), .D({ D[8:11] }), .ENP(N_6), .ENT(N_8),
            .LOAD(LOAD), .Q({ Q[8:11] }), .RCO(N_9) );
upflct4b QL4 ( .CLK(CLK), .CLR(CLR), .D({ D[4:7] }), .ENP(N_7), .ENT(N_10),
            .LOAD(LOAD), .Q({ Q[4:7] }), .RCO(N_8) );
upflct4c QL3 ( .CLK(CLK), .CLR(CLR), .D({ D[20:23] }), .ENP(N_1), .ENT(N_5),
            .LOAD(LOAD), .Q({ Q[20:23] }) );
upflcar2 QL2 ( .ACO1(N_7), .ACO2(N_6), .CLK(CLK), .CLR(CLR), .D({ D[0:1] }),
            .LOAD(LOAD) );
upflcar3 QL1 ( .ACO1(N_3), .ACO2(N_2), .ACO3(N_1), .CLK(CLK), .CLR(CLR),
            .D({ D[0:1] }), .LOAD(LOAD) );

endmodule // upflct24

`endif

`ifdef upflct16
`else
`define upflct16
module upflct16( CLK , CLR, D, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:15] D;
input LOAD;
 output [0:15] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;

upflct4a QL5 ( .CLK(CLK), .CLR(CLR), .D({ D[0:3] }), .LOAD(LOAD), .Q({ Q[0:3] }),
            .RCO(N_6) );
upflct4b QL4 ( .CLK(CLK), .CLR(CLR), .D({ D[8:11] }), .ENP(N_2), .ENT(N_4),
            .LOAD(LOAD), .Q({ Q[8:11] }), .RCO(N_5) );
upflct4b QL3 ( .CLK(CLK), .CLR(CLR), .D({ D[4:7] }), .ENP(N_3), .ENT(N_6),
            .LOAD(LOAD), .Q({ Q[4:7] }), .RCO(N_4) );
upflct4c QL2 ( .CLK(CLK), .CLR(CLR), .D({ D[12:15] }), .ENP(N_1), .ENT(N_5),
            .LOAD(LOAD), .Q({ Q[12:15] }) );
upflcar3 QL1 ( .ACO1(N_3), .ACO2(N_2), .ACO3(N_1), .CLK(CLK), .CLR(CLR),
            .D({ D[0:1] }), .LOAD(LOAD) );

endmodule // upflct16

`endif

`ifdef reg_lvpecl_outpad_25dc
`else
`define reg_lvpecl_outpad_25dc
module reg_lvpecl_outpad_25dc( clk , clr, input2diff, Vo_neg, Vo_pos );
input clk /* synthesis syn_isclock=1 */;
input clr /* synthesis syn_isclock=1 */;
input input2diff;
output Vo_neg, Vo_pos;
wire inv;
wire non_inv;
supply1 vcc;
supply0 gnd;

super_logic I4 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(gnd),
              .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd),
              .E1(gnd), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd),
              .F5(vcc), .F6(gnd), .MP(input2diff), .MS(gnd), .NP(input2diff),
              .NS(gnd), .NZ(inv), .OP(gnd), .OS(gnd), .OZ(non_inv), .PP(vcc),
              .PS(gnd), .QC(gnd), .QR(gnd), .QS(vcc) );
outpadff_25um I1 ( .A(inv), .FFCLK(clk), .FFCLR(clr), .P(Vo_neg) );
outpadff_25um I2 ( .A(non_inv), .FFCLK(clk), .FFCLR(clr), .P(Vo_pos) );

endmodule // reg_lvpecl_outpad_25dc

`endif

`ifdef reg_lvpecl_outpad_25ac
`else
`define reg_lvpecl_outpad_25ac
module reg_lvpecl_outpad_25ac( clk , clr, input2diff, Vo_neg, Vo_pos );
input input2diff;
input clk /* synthesis syn_isclock=1 */;
input clr /* synthesis syn_isclock=1 */;
output Vo_neg, Vo_pos;
wire inv;
wire non_inv;
supply1 vcc;
supply0 gnd;

eio_25um I8 ( .A2(gnd), .EN(vcc), .FFCLK(clk), .FFCLR(clr), .I_EN(gnd),
           .OE_EN(non_inv), .OESEL(gnd), .OSEL(vcc), .P(Vo_neg) );
eio_25um I9 ( .A2(gnd), .EN(vcc), .FFCLK(clk), .FFCLR(clr), .I_EN(gnd),
           .OE_EN(inv), .OESEL(gnd), .OSEL(vcc), .P(Vo_pos) );
super_logic I4 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(gnd),
              .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd),
              .E1(gnd), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd),
              .F5(vcc), .F6(gnd), .MP(input2diff), .MS(gnd), .NP(input2diff),
              .NS(gnd), .NZ(inv), .OP(gnd), .OS(gnd), .OZ(non_inv), .PP(vcc),
              .PS(gnd), .QC(gnd), .QR(gnd), .QS(vcc) );

endmodule // reg_lvpecl_outpad_25ac

`endif

`ifdef lvpecl_outpad_25dc
`else
`define lvpecl_outpad_25dc
module lvpecl_outpad_25dc( input2diff , Vo_neg, Vo_pos );
input input2diff;
output Vo_neg, Vo_pos;
wire inv;
wire non_inv;
supply1 vcc;
supply0 gnd;

outpad_25um I5 ( .A(inv), .P(Vo_neg) );
outpad_25um I6 ( .A(non_inv), .P(Vo_pos) );
super_logic I4 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(gnd),
              .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd),
              .E1(gnd), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd),
              .F5(vcc), .F6(gnd), .MP(input2diff), .MS(gnd), .NP(input2diff),
              .NS(gnd), .NZ(inv), .OP(gnd), .OS(gnd), .OZ(non_inv), .PP(vcc),
              .PS(gnd), .QC(gnd), .QR(gnd), .QS(vcc) );

endmodule // lvpecl_outpad_25dc

`endif

`ifdef lvpecl_outpad_25ac
`else
`define lvpecl_outpad_25ac
module lvpecl_outpad_25ac( input2diff , Vo_neg, Vo_pos );
input input2diff;
output Vo_neg, Vo_pos;
wire inv;
wire non_inv;
supply1 vcc;
supply0 gnd;

tripadod_25um I7 ( .EN(non_inv), .P(Vo_neg) );
tripadod_25um I8 ( .EN(inv), .P(Vo_pos) );
super_logic I9 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(gnd),
              .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd),
              .E1(gnd), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd),
              .F5(vcc), .F6(gnd), .MP(input2diff), .MS(gnd), .NP(input2diff),
              .NS(gnd), .NZ(inv), .OP(gnd), .OS(gnd), .OZ(non_inv), .PP(vcc),
              .PS(gnd), .QC(gnd), .QR(gnd), .QS(vcc) );

endmodule // lvpecl_outpad_25ac

`endif

`ifdef lvpecl_inpad_25
`else
`define lvpecl_inpad_25
module lvpecl_inpad_25( Vin_neg , Vin_pos, diff_input );
output diff_input;
input Vin_neg, Vin_pos;
wire N_1;
wire N_2;

and2i1 I5 ( .A(N_1), .B(N_2), .Q(diff_input) );
inpad_25um I6 ( .P(Vin_neg), .Q(N_2) );
inpad_25um I7 ( .P(Vin_pos), .Q(N_1) );

endmodule // lvpecl_inpad_25

`endif

`ifdef reg_lvds_outpad_25dc
`else
`define reg_lvds_outpad_25dc
module reg_lvds_outpad_25dc( clk , clr, input2diff, Vo_neg, Vo_pos );
input clk /* synthesis syn_isclock=1 */;
input clr /* synthesis syn_isclock=1 */;
input input2diff;
output Vo_neg, Vo_pos;
wire inv;
wire non_inv;
supply1 vcc;
supply0 gnd;

super_logic I4 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(gnd),
              .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd),
              .E1(gnd), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd),
              .F5(vcc), .F6(gnd), .MP(input2diff), .MS(gnd), .NP(input2diff),
              .NS(gnd), .NZ(inv), .OP(gnd), .OS(gnd), .OZ(non_inv), .PP(vcc),
              .PS(gnd), .QC(gnd), .QR(gnd), .QS(vcc) );
outpadff_25um I2 ( .A(non_inv), .FFCLK(clk), .FFCLR(clr), .P(Vo_pos) );
outpadff_25um I1 ( .A(inv), .FFCLK(clk), .FFCLR(clr), .P(Vo_neg) );

endmodule // reg_lvds_outpad_25dc

`endif

`ifdef lvds_outpad_25dc
`else
`define lvds_outpad_25dc
module lvds_outpad_25dc( input2diff , Vo_neg, Vo_pos );
input input2diff;
output Vo_neg, Vo_pos;
wire inv;
wire non_inv;
supply1 vcc;
supply0 gnd;

outpad_25um I5 ( .A(inv), .P(Vo_neg) );
outpad_25um I6 ( .A(non_inv), .P(Vo_pos) );
super_logic I4 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(gnd),
              .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd),
              .E1(gnd), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd),
              .F5(vcc), .F6(gnd), .MP(input2diff), .MS(gnd), .NP(input2diff),
              .NS(gnd), .NZ(inv), .OP(gnd), .OS(gnd), .OZ(non_inv), .PP(vcc),
              .PS(gnd), .QC(gnd), .QR(gnd), .QS(vcc) );

endmodule // lvds_outpad_25dc

`endif

`ifdef lvds_inpad_25dc
`else
`define lvds_inpad_25dc
module lvds_inpad_25dc( Vin_neg , Vin_pos, diff_input );
output diff_input;
input Vin_neg, Vin_pos;
wire N_1;
wire N_2;

and2i1 I5 ( .A(N_1), .B(N_2), .Q(diff_input) );
inpad_25um I6 ( .P(Vin_neg), .Q(N_2) );
inpad_25um I7 ( .P(Vin_pos), .Q(N_1) );

endmodule // lvds_inpad_25dc

`endif

`ifdef uct8p2
`else
`define uct8p2
module uct8p2( CLK , CLR, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 output [7:0] Q;
wire Q1Q2Q3;
wire N_1;
supply0 GND;
wire UCTCO;
supply1 VCC;

mux2x2 I_60 ( .A(GND), .B(Q[0]), .Q(N_1), .S(Q1Q2Q3) );
dffc I_61 ( .CLK(CLK), .CLR(CLR), .D(N_1), .Q(UCTCO) );
and3i0 I_17 ( .A(Q[1]), .B(Q[2]), .C(Q[3]), .Q(Q1Q2Q3) );
ucebit2a UCT4 ( .CLK(CLK), .CLR(CLR), .ENH1(UCTCO), .ENH2(VCC), .ENH3(VCC),
             .ENH4(VCC), .ENL1(GND), .ENL2(GND), .ENL3(GND), .Q(Q[4]),
             .QFB(Q[4]) );
ucebit2a UCT0 ( .CLK(CLK), .CLR(CLR), .ENH1(VCC), .ENH2(VCC), .ENH3(VCC),
             .ENH4(VCC), .ENL1(GND), .ENL2(GND), .ENL3(GND), .Q(Q[0]),
             .QFB(Q[0]) );
ucebit2a UCT7 ( .CLK(CLK), .CLR(CLR), .ENH1(Q[4]), .ENH2(Q[5]), .ENH3(Q[6]),
             .ENH4(UCTCO), .ENL1(GND), .ENL2(GND), .ENL3(GND), .Q(Q[7]),
             .QFB(Q[7]) );
ucebit2a UCT6 ( .CLK(CLK), .CLR(CLR), .ENH1(Q[4]), .ENH2(Q[5]), .ENH3(UCTCO),
             .ENH4(VCC), .ENL1(GND), .ENL2(GND), .ENL3(GND), .Q(Q[6]),
             .QFB(Q[6]) );
ucebit2a UCT5 ( .CLK(CLK), .CLR(CLR), .ENH1(Q[4]), .ENH2(UCTCO), .ENH3(VCC),
             .ENH4(VCC), .ENL1(GND), .ENL2(GND), .ENL3(GND), .Q(Q[5]),
             .QFB(Q[5]) );
ucebit2a UCT3 ( .CLK(CLK), .CLR(CLR), .ENH1(Q[0]), .ENH2(Q[1]), .ENH3(Q[2]),
             .ENH4(VCC), .ENL1(GND), .ENL2(GND), .ENL3(GND), .Q(Q[3]),
             .QFB(Q[3]) );
ucebit2a UCT2 ( .CLK(CLK), .CLR(CLR), .ENH1(Q[0]), .ENH2(Q[1]), .ENH3(VCC),
             .ENH4(VCC), .ENL1(GND), .ENL2(GND), .ENL3(GND), .Q(Q[2]),
             .QFB(Q[2]) );
ucebit2a UCT1 ( .CLK(CLK), .CLR(CLR), .ENH1(Q[0]), .ENH2(VCC), .ENH3(VCC),
             .ENH4(VCC), .ENL1(GND), .ENL2(GND), .ENL3(GND), .Q(Q[1]),
             .QFB(Q[1]) );

endmodule // uct8p2

`endif

`ifdef tpad8_25um
`else
`define tpad8_25um
module tpad8_25um( A , EN, P );
 input [7:0] A;
input EN;
 output [7:0] P;

tripad_25um I1 ( .A(A[0]), .EN(EN), .P(P[0]) );
tripad_25um I2 ( .A(A[1]), .EN(EN), .P(P[1]) );
tripad_25um I3 ( .A(A[2]), .EN(EN), .P(P[2]) );
tripad_25um I4 ( .A(A[3]), .EN(EN), .P(P[3]) );
tripad_25um I5 ( .A(A[4]), .EN(EN), .P(P[4]) );
tripad_25um I6 ( .A(A[5]), .EN(EN), .P(P[5]) );
tripad_25um I7 ( .A(A[6]), .EN(EN), .P(P[6]) );
tripad_25um I8 ( .A(A[7]), .EN(EN), .P(P[7]) );

endmodule // tpad8_25um

`endif

`ifdef tpad8ff_25um
`else
`define tpad8ff_25um
module tpad8ff_25um( A , EN, FFCLK, FFCLR, P, Q );
 input [7:0] A;
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input EN;
 output [7:0] P;
 output [7:0] Q;

tripadff_25um I4 ( .A(A[3]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[3]),
                .Q(Q[3]) );
tripadff_25um I3 ( .A(A[2]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[2]),
                .Q(Q[2]) );
tripadff_25um I2 ( .A(A[1]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[1]),
                .Q(Q[1]) );
tripadff_25um I1 ( .A(A[0]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[0]),
                .Q(Q[0]) );
tripadff_25um I5 ( .A(A[4]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[4]),
                .Q(Q[4]) );
tripadff_25um I6 ( .A(A[5]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[5]),
                .Q(Q[5]) );
tripadff_25um I7 ( .A(A[6]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[6]),
                .Q(Q[6]) );
tripadff_25um I8 ( .A(A[7]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[7]),
                .Q(Q[7]) );

endmodule // tpad8ff_25um

`endif

`ifdef tpad4ff_25um
`else
`define tpad4ff_25um
module tpad4ff_25um( A , EN, FFCLK, FFCLR, P, Q );
 input [3:0] A;
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input EN;
 output [3:0] P;
 output [3:0] Q;

tripadff_25um I1 ( .A(A[0]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[0]),
                .Q(Q[0]) );
tripadff_25um I2 ( .A(A[1]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[1]),
                .Q(Q[1]) );
tripadff_25um I3 ( .A(A[2]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[2]),
                .Q(Q[2]) );
tripadff_25um I4 ( .A(A[3]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[3]),
                .Q(Q[3]) );

endmodule // tpad4ff_25um

`endif

`ifdef tpad4_25um
`else
`define tpad4_25um
module tpad4_25um( A , EN, P );
 input [3:0] A;
input EN;
 output [3:0] P;

tripad_25um I1 ( .A(A[0]), .EN(EN), .P(P[0]) );
tripad_25um I2 ( .A(A[1]), .EN(EN), .P(P[1]) );
tripad_25um I3 ( .A(A[2]), .EN(EN), .P(P[2]) );
tripad_25um I4 ( .A(A[3]), .EN(EN), .P(P[3]) );

endmodule // tpad4_25um

`endif

`ifdef tpad16ff_25um
`else
`define tpad16ff_25um
module tpad16ff_25um( A , EN, FFCLK, FFCLR, P, Q );
 input [15:0] A;
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input EN;
 output [15:0] P;
 output [15:0] Q;

tripadff_25um I1 ( .A(A[0]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[0]),
                .Q(Q[0]) );
tripadff_25um I2 ( .A(A[1]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[1]),
                .Q(Q[1]) );
tripadff_25um I3 ( .A(A[2]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[2]),
                .Q(Q[2]) );
tripadff_25um I10 ( .A(A[3]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[3]),
                 .Q(Q[3]) );
tripadff_25um I4 ( .A(A[4]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[4]),
                .Q(Q[4]) );
tripadff_25um I5 ( .A(A[5]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[5]),
                .Q(Q[5]) );
tripadff_25um I6 ( .A(A[6]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[6]),
                .Q(Q[6]) );
tripadff_25um I11 ( .A(A[7]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[7]),
                 .Q(Q[7]) );
tripadff_25um I7 ( .A(A[8]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[8]),
                .Q(Q[8]) );
tripadff_25um I8 ( .A(A[9]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[9]),
                .Q(Q[9]) );
tripadff_25um I9 ( .A(A[10]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[10]),
                .Q(Q[10]) );
tripadff_25um I12 ( .A(A[11]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[11]),
                 .Q(Q[11]) );
tripadff_25um I13 ( .A(A[12]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[12]),
                 .Q(Q[12]) );
tripadff_25um I14 ( .A(A[13]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[13]),
                 .Q(Q[13]) );
tripadff_25um I15 ( .A(A[14]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[14]),
                 .Q(Q[14]) );
tripadff_25um I16 ( .A(A[15]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[15]),
                 .Q(Q[15]) );

endmodule // tpad16ff_25um

`endif

`ifdef tpad16_25um
`else
`define tpad16_25um
module tpad16_25um( A , EN, P );
 input [15:0] A;
input EN;
 output [15:0] P;

tripad_25um I1 ( .A(A[0]), .EN(EN), .P(P[0]) );
tripad_25um I2 ( .A(A[1]), .EN(EN), .P(P[1]) );
tripad_25um I3 ( .A(A[2]), .EN(EN), .P(P[2]) );
tripad_25um I4 ( .A(A[3]), .EN(EN), .P(P[3]) );
tripad_25um I5 ( .A(A[4]), .EN(EN), .P(P[4]) );
tripad_25um I6 ( .A(A[5]), .EN(EN), .P(P[5]) );
tripad_25um I7 ( .A(A[6]), .EN(EN), .P(P[6]) );
tripad_25um I8 ( .A(A[7]), .EN(EN), .P(P[7]) );
tripad_25um I9 ( .A(A[8]), .EN(EN), .P(P[8]) );
tripad_25um I10 ( .A(A[9]), .EN(EN), .P(P[9]) );
tripad_25um I11 ( .A(A[10]), .EN(EN), .P(P[10]) );
tripad_25um I12 ( .A(A[11]), .EN(EN), .P(P[11]) );
tripad_25um I13 ( .A(A[12]), .EN(EN), .P(P[12]) );
tripad_25um I14 ( .A(A[13]), .EN(EN), .P(P[13]) );
tripad_25um I15 ( .A(A[14]), .EN(EN), .P(P[14]) );
tripad_25um I16 ( .A(A[15]), .EN(EN), .P(P[15]) );

endmodule // tpad16_25um

`endif

`ifdef opad8ff_25um
`else
`define opad8ff_25um
module opad8ff_25um( A , FFCLK, FFCLR, P, P_FB );
 input [7:0] A;
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
 output [7:0] P;
 output [7:0] P_FB;

outpadff_25um I1 ( .A(A[0]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[0]),
                .P_FB(P_FB[0]) );
outpadff_25um I2 ( .A(A[1]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[1]),
                .P_FB(P_FB[1]) );
outpadff_25um I3 ( .A(A[2]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[2]),
                .P_FB(P_FB[2]) );
outpadff_25um I4 ( .A(A[3]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[3]),
                .P_FB(P_FB[3]) );
outpadff_25um I5 ( .A(A[4]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[4]),
                .P_FB(P_FB[4]) );
outpadff_25um I6 ( .A(A[5]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[5]),
                .P_FB(P_FB[5]) );
outpadff_25um I7 ( .A(A[6]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[6]),
                .P_FB(P_FB[6]) );
outpadff_25um I8 ( .A(A[7]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[7]),
                .P_FB(P_FB[7]) );

endmodule // opad8ff_25um

`endif

`ifdef opad8_25um
`else
`define opad8_25um
module opad8_25um( A , P );
 input [7:0] A;
 output [7:0] P;

outpad_25um I1 ( .A(A[0]), .P(P[0]) );
outpad_25um I2 ( .A(A[1]), .P(P[1]) );
outpad_25um I3 ( .A(A[2]), .P(P[2]) );
outpad_25um I4 ( .A(A[3]), .P(P[3]) );
outpad_25um I5 ( .A(A[4]), .P(P[4]) );
outpad_25um I6 ( .A(A[5]), .P(P[5]) );
outpad_25um I7 ( .A(A[6]), .P(P[6]) );
outpad_25um I8 ( .A(A[7]), .P(P[7]) );

endmodule // opad8_25um

`endif

`ifdef opad4ff_25um
`else
`define opad4ff_25um
module opad4ff_25um( A , FFCLK, FFCLR, P, P_FB );
 input [3:0] A;
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
 output [3:0] P;
 output [3:0] P_FB;

outpadff_25um I1 ( .A(A[0]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[0]),
                .P_FB(P_FB[0]) );
outpadff_25um I2 ( .A(A[1]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[1]),
                .P_FB(P_FB[1]) );
outpadff_25um I3 ( .A(A[2]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[2]),
                .P_FB(P_FB[2]) );
outpadff_25um I4 ( .A(A[3]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[3]),
                .P_FB(P_FB[3]) );

endmodule // opad4ff_25um

`endif

`ifdef opad4_25um
`else
`define opad4_25um
module opad4_25um( A , P );
 input [3:0] A;
 output [3:0] P;

outpad_25um I1 ( .A(A[0]), .P(P[0]) );
outpad_25um I2 ( .A(A[1]), .P(P[1]) );
outpad_25um I3 ( .A(A[2]), .P(P[2]) );
outpad_25um I4 ( .A(A[3]), .P(P[3]) );

endmodule // opad4_25um

`endif

`ifdef opad16ff_25um
`else
`define opad16ff_25um
module opad16ff_25um( A , FFCLK, FFCLR, P, P_FB );
 input [15:0] A;
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
 output [15:0] P;
 output [15:0] P_FB;

outpadff_25um I4 ( .A(A[0]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[0]),
                .P_FB(P_FB[0]) );
outpadff_25um I1 ( .A(A[1]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[1]),
                .P_FB(P_FB[1]) );
outpadff_25um I2 ( .A(A[2]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[2]),
                .P_FB(P_FB[2]) );
outpadff_25um I3 ( .A(A[3]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[3]),
                .P_FB(P_FB[3]) );
outpadff_25um I5 ( .A(A[4]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[4]),
                .P_FB(P_FB[4]) );
outpadff_25um I6 ( .A(A[5]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[5]),
                .P_FB(P_FB[5]) );
outpadff_25um I7 ( .A(A[6]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[6]),
                .P_FB(P_FB[6]) );
outpadff_25um I8 ( .A(A[7]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[7]),
                .P_FB(P_FB[7]) );
outpadff_25um I13 ( .A(A[8]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[8]),
                 .P_FB(P_FB[8]) );
outpadff_25um I14 ( .A(A[9]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[9]),
                 .P_FB(P_FB[9]) );
outpadff_25um I15 ( .A(A[10]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[10]),
                 .P_FB(P_FB[10]) );
outpadff_25um I16 ( .A(A[11]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[11]),
                 .P_FB(P_FB[11]) );
outpadff_25um I9 ( .A(A[12]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[12]),
                .P_FB(P_FB[12]) );
outpadff_25um I10 ( .A(A[13]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[13]),
                 .P_FB(P_FB[13]) );
outpadff_25um I11 ( .A(A[14]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[14]),
                 .P_FB(P_FB[14]) );
outpadff_25um I12 ( .A(A[15]), .FFCLK(FFCLK), .FFCLR(FFCLR), .P(P[15]),
                 .P_FB(P_FB[15]) );

endmodule // opad16ff_25um

`endif

`ifdef opad16_25um
`else
`define opad16_25um
module opad16_25um( A , P );
 input [15:0] A;
 output [15:0] P;

outpad_25um I1 ( .A(A[0]), .P(P[0]) );
outpad_25um I2 ( .A(A[1]), .P(P[1]) );
outpad_25um I3 ( .A(A[2]), .P(P[2]) );
outpad_25um I4 ( .A(A[3]), .P(P[3]) );
outpad_25um I5 ( .A(A[4]), .P(P[4]) );
outpad_25um I6 ( .A(A[5]), .P(P[5]) );
outpad_25um I7 ( .A(A[6]), .P(P[6]) );
outpad_25um I8 ( .A(A[7]), .P(P[7]) );
outpad_25um I9 ( .A(A[8]), .P(P[8]) );
outpad_25um I10 ( .A(A[9]), .P(P[9]) );
outpad_25um I11 ( .A(A[10]), .P(P[10]) );
outpad_25um I12 ( .A(A[11]), .P(P[11]) );
outpad_25um I13 ( .A(A[12]), .P(P[12]) );
outpad_25um I14 ( .A(A[13]), .P(P[13]) );
outpad_25um I15 ( .A(A[14]), .P(P[14]) );
outpad_25um I16 ( .A(A[15]), .P(P[15]) );

endmodule // opad16_25um

`endif

`ifdef ipad8ff_25um
`else
`define ipad8ff_25um
module ipad8ff_25um( FFCLK , FFCLR, FFEN, P, FFQ, Q );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input FFEN;
 output [7:0] FFQ;
 input [7:0] P;
 output [7:0] Q;

inpadff_25um I7 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[0]),
               .P(P[0]), .Q(Q[0]) );
inpadff_25um I6 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[1]),
               .P(P[1]), .Q(Q[1]) );
inpadff_25um I5 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[2]),
               .P(P[2]), .Q(Q[2]) );
inpadff_25um I4 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[3]),
               .P(P[3]), .Q(Q[3]) );
inpadff_25um I8 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[4]),
               .P(P[4]), .Q(Q[4]) );
inpadff_25um I9 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[5]),
               .P(P[5]), .Q(Q[5]) );
inpadff_25um I10 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[6]),
                .P(P[6]), .Q(Q[6]) );
inpadff_25um I11 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[7]),
                .P(P[7]), .Q(Q[7]) );

endmodule // ipad8ff_25um

`endif

`ifdef ipad8_25um
`else
`define ipad8_25um
module ipad8_25um( P , Q );
 input [7:0] P;
 output [7:0] Q;

inpad_25um I1 ( .P(P[4]), .Q(Q[4]) );
inpad_25um I2 ( .P(P[5]), .Q(Q[5]) );
inpad_25um I3 ( .P(P[6]), .Q(Q[6]) );
inpad_25um I4 ( .P(P[7]), .Q(Q[7]) );
inpad_25um I5 ( .P(P[3]), .Q(Q[3]) );
inpad_25um I6 ( .P(P[2]), .Q(Q[2]) );
inpad_25um I7 ( .P(P[1]), .Q(Q[1]) );
inpad_25um I8 ( .P(P[0]), .Q(Q[0]) );

endmodule // ipad8_25um

`endif

`ifdef ipad4ff_25um
`else
`define ipad4ff_25um
module ipad4ff_25um( FFCLK , FFCLR, FFEN, P, FFQ, Q );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input FFEN;
 output [3:0] FFQ;
 input [3:0] P;
 output [3:0] Q;

inpadff_25um I4 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[3]),
               .P(P[3]), .Q(Q[3]) );
inpadff_25um I1 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[0]),
               .P(P[0]), .Q(Q[0]) );
inpadff_25um I2 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[1]),
               .P(P[1]), .Q(Q[1]) );
inpadff_25um I3 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[2]),
               .P(P[2]), .Q(Q[2]) );

endmodule // ipad4ff_25um

`endif

`ifdef ipad4_25um
`else
`define ipad4_25um
module ipad4_25um( P , Q );
 input [3:0] P;
 output [3:0] Q;

inpad_25um I1 ( .P(P[3]), .Q(Q[3]) );
inpad_25um I2 ( .P(P[2]), .Q(Q[2]) );
inpad_25um I3 ( .P(P[1]), .Q(Q[1]) );
inpad_25um I4 ( .P(P[0]), .Q(Q[0]) );

endmodule // ipad4_25um

`endif

`ifdef ipad16ff_25um
`else
`define ipad16ff_25um
module ipad16ff_25um( FFCLK , FFCLR, FFEN, P, FFQ, Q );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input FFEN;
 output [15:0] FFQ;
 input [15:0] P;
 output [15:0] Q;

inpadff_25um I9 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[0]),
               .P(P[0]), .Q(Q[0]) );
inpadff_25um I10 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[1]),
                .P(P[1]), .Q(Q[1]) );
inpadff_25um I11 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[2]),
                .P(P[2]), .Q(Q[2]) );
inpadff_25um I12 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[3]),
                .P(P[3]), .Q(Q[3]) );
inpadff_25um I13 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[4]),
                .P(P[4]), .Q(Q[4]) );
inpadff_25um I14 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[5]),
                .P(P[5]), .Q(Q[5]) );
inpadff_25um I15 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[6]),
                .P(P[6]), .Q(Q[6]) );
inpadff_25um I16 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[7]),
                .P(P[7]), .Q(Q[7]) );
inpadff_25um I17 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[8]),
                .P(P[8]), .Q(Q[8]) );
inpadff_25um I18 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[9]),
                .P(P[9]), .Q(Q[9]) );
inpadff_25um I19 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[10]),
                .P(P[10]), .Q(Q[10]) );
inpadff_25um I20 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[11]),
                .P(P[11]), .Q(Q[11]) );
inpadff_25um I21 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[12]),
                .P(P[12]), .Q(Q[12]) );
inpadff_25um I22 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[13]),
                .P(P[13]), .Q(Q[13]) );
inpadff_25um I23 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[14]),
                .P(P[14]), .Q(Q[14]) );
inpadff_25um I24 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[15]),
                .P(P[15]), .Q(Q[15]) );

endmodule // ipad16ff_25um

`endif

`ifdef ipad16_25um
`else
`define ipad16_25um
module ipad16_25um( P , Q );
 input [15:0] P;
 output [15:0] Q;

inpad_25um I1 ( .P(P[15]), .Q(Q[15]) );
inpad_25um I2 ( .P(P[14]), .Q(Q[14]) );
inpad_25um I3 ( .P(P[13]), .Q(Q[13]) );
inpad_25um I4 ( .P(P[12]), .Q(Q[12]) );
inpad_25um I5 ( .P(P[8]), .Q(Q[8]) );
inpad_25um I6 ( .P(P[9]), .Q(Q[9]) );
inpad_25um I7 ( .P(P[10]), .Q(Q[10]) );
inpad_25um I8 ( .P(P[11]), .Q(Q[11]) );
inpad_25um I9 ( .P(P[7]), .Q(Q[7]) );
inpad_25um I10 ( .P(P[6]), .Q(Q[6]) );
inpad_25um I11 ( .P(P[5]), .Q(Q[5]) );
inpad_25um I12 ( .P(P[4]), .Q(Q[4]) );
inpad_25um I13 ( .P(P[3]), .Q(Q[3]) );
inpad_25um I14 ( .P(P[2]), .Q(Q[2]) );
inpad_25um I15 ( .P(P[1]), .Q(Q[1]) );
inpad_25um I16 ( .P(P[0]), .Q(Q[0]) );

endmodule // ipad16_25um

`endif

`ifdef bpad8iff_25um
`else
`define bpad8iff_25um
module bpad8iff_25um( A2 , EN, FFCLK, FFCLR, FFEN, FFQ, Q, P );
 input [7:0] A2;
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input EN, FFEN;
 output [7:0] FFQ;
 inout [7:0] P;
 output [7:0] Q;

bipadiff_25um I24 ( .A2(A2[0]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[0]), .P(P[0]), .Q(Q[0]) );
bipadiff_25um I25 ( .A2(A2[1]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[1]), .P(P[1]), .Q(Q[1]) );
bipadiff_25um I26 ( .A2(A2[2]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[2]), .P(P[2]), .Q(Q[2]) );
bipadiff_25um I27 ( .A2(A2[3]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[3]), .P(P[3]), .Q(Q[3]) );
bipadiff_25um I28 ( .A2(A2[4]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[4]), .P(P[4]), .Q(Q[4]) );
bipadiff_25um I29 ( .A2(A2[5]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[5]), .P(P[5]), .Q(Q[5]) );
bipadiff_25um I30 ( .A2(A2[6]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[6]), .P(P[6]), .Q(Q[6]) );
bipadiff_25um I31 ( .A2(A2[7]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[7]), .P(P[7]), .Q(Q[7]) );

endmodule // bpad8iff_25um

`endif

`ifdef bpad8_25um
`else
`define bpad8_25um
module bpad8_25um( A , EN, Q, P );
 input [7:0] A;
input EN;
 inout [7:0] P;
 output [7:0] Q;

bipad_25um I1 ( .A(A[4]), .EN(EN), .P(P[4]), .Q(Q[4]) );
bipad_25um I2 ( .A(A[5]), .EN(EN), .P(P[5]), .Q(Q[5]) );
bipad_25um I3 ( .A(A[6]), .EN(EN), .P(P[6]), .Q(Q[6]) );
bipad_25um I4 ( .A(A[7]), .EN(EN), .P(P[7]), .Q(Q[7]) );
bipad_25um I5 ( .A(A[3]), .EN(EN), .P(P[3]), .Q(Q[3]) );
bipad_25um I6 ( .A(A[2]), .EN(EN), .P(P[2]), .Q(Q[2]) );
bipad_25um I7 ( .A(A[1]), .EN(EN), .P(P[1]), .Q(Q[1]) );
bipad_25um I8 ( .A(A[0]), .EN(EN), .P(P[0]), .Q(Q[0]) );

endmodule // bpad8_25um

`endif

`ifdef bpad4iff_25um
`else
`define bpad4iff_25um
module bpad4iff_25um( A2 , EN, FFCLK, FFCLR, FFEN, FFQ, Q, P );
 input [3:0] A2;
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input EN, FFEN;
 output [3:0] FFQ;
 inout [3:0] P;
 output [3:0] Q;

bipadiff_25um I18 ( .A2(A2[0]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[0]), .P(P[0]), .Q(Q[0]) );
bipadiff_25um I19 ( .A2(A2[1]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[1]), .P(P[1]), .Q(Q[1]) );
bipadiff_25um I20 ( .A2(A2[2]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[2]), .P(P[2]), .Q(Q[2]) );
bipadiff_25um I21 ( .A2(A2[3]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[3]), .P(P[3]), .Q(Q[3]) );

endmodule // bpad4iff_25um

`endif

`ifdef bpad4_25um
`else
`define bpad4_25um
module bpad4_25um( A , EN, Q, P );
 input [3:0] A;
input EN;
 inout [3:0] P;
 output [3:0] Q;

bipad_25um I1 ( .A(A[3]), .EN(EN), .P(P[3]), .Q(Q[3]) );
bipad_25um I2 ( .A(A[2]), .EN(EN), .P(P[2]), .Q(Q[2]) );
bipad_25um I3 ( .A(A[1]), .EN(EN), .P(P[1]), .Q(Q[1]) );
bipad_25um I4 ( .A(A[0]), .EN(EN), .P(P[0]), .Q(Q[0]) );

endmodule // bpad4_25um

`endif

`ifdef bpad16iff_25um
`else
`define bpad16iff_25um
module bpad16iff_25um( A2 , EN, FFCLK, FFCLR, FFEN, FFQ, Q, P );
 input [15:0] A2;
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input EN, FFEN;
 output [15:0] FFQ;
 inout [15:0] P;
 output [15:0] Q;

bipadiff_25um I39 ( .A2(A2[0]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[0]), .P(P[0]), .Q(Q[0]) );
bipadiff_25um I38 ( .A2(A2[1]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[1]), .P(P[1]), .Q(Q[1]) );
bipadiff_25um I37 ( .A2(A2[2]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[2]), .P(P[2]), .Q(Q[2]) );
bipadiff_25um I36 ( .A2(A2[3]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[3]), .P(P[3]), .Q(Q[3]) );
bipadiff_25um I40 ( .A2(A2[4]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[4]), .P(P[4]), .Q(Q[4]) );
bipadiff_25um I41 ( .A2(A2[5]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[5]), .P(P[5]), .Q(Q[5]) );
bipadiff_25um I42 ( .A2(A2[6]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[6]), .P(P[6]), .Q(Q[6]) );
bipadiff_25um I43 ( .A2(A2[7]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[7]), .P(P[7]), .Q(Q[7]) );
bipadiff_25um I47 ( .A2(A2[8]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[8]), .P(P[8]), .Q(Q[8]) );
bipadiff_25um I46 ( .A2(A2[9]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[9]), .P(P[9]), .Q(Q[9]) );
bipadiff_25um I45 ( .A2(A2[10]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[10]), .P(P[10]), .Q(Q[10]) );
bipadiff_25um I44 ( .A2(A2[11]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[11]), .P(P[11]), .Q(Q[11]) );
bipadiff_25um I48 ( .A2(A2[12]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[12]), .P(P[12]), .Q(Q[12]) );
bipadiff_25um I49 ( .A2(A2[13]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[13]), .P(P[13]), .Q(Q[13]) );
bipadiff_25um I50 ( .A2(A2[14]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[14]), .P(P[14]), .Q(Q[14]) );
bipadiff_25um I51 ( .A2(A2[15]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR),
                 .FFEN(FFEN), .FFQ(FFQ[15]), .P(P[15]), .Q(Q[15]) );

endmodule // bpad16iff_25um

`endif

`ifdef bpad16_25um
`else
`define bpad16_25um
module bpad16_25um( A , EN, Q, P );
 input [15:0] A;
input EN;
 inout [15:0] P;
 output [15:0] Q;

bipad_25um I1 ( .A(A[12]), .EN(EN), .P(P[12]), .Q(Q[12]) );
bipad_25um I2 ( .A(A[13]), .EN(EN), .P(P[13]), .Q(Q[13]) );
bipad_25um I3 ( .A(A[14]), .EN(EN), .P(P[14]), .Q(Q[14]) );
bipad_25um I4 ( .A(A[15]), .EN(EN), .P(P[15]), .Q(Q[15]) );
bipad_25um I5 ( .A(A[11]), .EN(EN), .P(P[11]), .Q(Q[11]) );
bipad_25um I6 ( .A(A[10]), .EN(EN), .P(P[10]), .Q(Q[10]) );
bipad_25um I7 ( .A(A[9]), .EN(EN), .P(P[9]), .Q(Q[9]) );
bipad_25um I8 ( .A(A[8]), .EN(EN), .P(P[8]), .Q(Q[8]) );
bipad_25um I9 ( .A(A[4]), .EN(EN), .P(P[4]), .Q(Q[4]) );
bipad_25um I10 ( .A(A[5]), .EN(EN), .P(P[5]), .Q(Q[5]) );
bipad_25um I11 ( .A(A[6]), .EN(EN), .P(P[6]), .Q(Q[6]) );
bipad_25um I12 ( .A(A[7]), .EN(EN), .P(P[7]), .Q(Q[7]) );
bipad_25um I13 ( .A(A[3]), .EN(EN), .P(P[3]), .Q(Q[3]) );
bipad_25um I14 ( .A(A[2]), .EN(EN), .P(P[2]), .Q(Q[2]) );
bipad_25um I15 ( .A(A[1]), .EN(EN), .P(P[1]), .Q(Q[1]) );
bipad_25um I16 ( .A(A[0]), .EN(EN), .P(P[0]), .Q(Q[0]) );

endmodule // bpad16_25um

`endif

`ifdef rgec8_25um
`else
`define rgec8_25um
module rgec8_25um( CLK , CLR, D, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [7:0] D;
input EN;
 output [7:0] Q;
supply0 gnd;

dffepc_2 I6 ( .CLK(CLK), .CLR(CLR), .D1(D[6]), .D2(D[7]), .EN1(EN), .EN2(EN),
           .PRE(gnd), .Q1(Q[6]), .Q2(Q[7]) );
dffepc_2 I7 ( .CLK(CLK), .CLR(CLR), .D1(D[4]), .D2(D[5]), .EN1(EN), .EN2(EN),
           .PRE(gnd), .Q1(Q[4]), .Q2(Q[5]) );
dffepc_2 I8 ( .CLK(CLK), .CLR(CLR), .D1(D[2]), .D2(D[3]), .EN1(EN), .EN2(EN),
           .PRE(gnd), .Q1(Q[2]), .Q2(Q[3]) );
dffepc_2 I9 ( .CLK(CLK), .CLR(CLR), .D1(D[0]), .D2(D[1]), .EN1(EN), .EN2(EN),
           .PRE(gnd), .Q1(Q[0]), .Q2(Q[1]) );

endmodule // rgec8_25um

`endif

`ifdef rgec4_25um
`else
`define rgec4_25um
module rgec4_25um( CLK , CLR, D, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [3:0] D;
input EN;
 output [3:0] Q;
supply0 gnd;

dffepc_2 I8 ( .CLK(CLK), .CLR(CLR), .D1(D[2]), .D2(D[3]), .EN1(EN), .EN2(EN),
           .PRE(gnd), .Q1(Q[2]), .Q2(Q[3]) );
dffepc_2 I9 ( .CLK(CLK), .CLR(CLR), .D1(D[0]), .D2(D[1]), .EN1(EN), .EN2(EN),
           .PRE(gnd), .Q1(Q[0]), .Q2(Q[1]) );

endmodule // rgec4_25um

`endif

`ifdef rgec16_25um
`else
`define rgec16_25um
module rgec16_25um( CLK , CLR, D, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [15:0] D;
input EN;
 output [15:0] Q;
supply0 gnd;

dffepc_2 I2 ( .CLK(CLK), .CLR(CLR), .D1(D[14]), .D2(D[15]), .EN1(EN), .EN2(EN),
           .PRE(gnd), .Q1(Q[14]), .Q2(Q[15]) );
dffepc_2 I3 ( .CLK(CLK), .CLR(CLR), .D1(D[12]), .D2(D[13]), .EN1(EN), .EN2(EN),
           .PRE(gnd), .Q1(Q[12]), .Q2(Q[13]) );
dffepc_2 I4 ( .CLK(CLK), .CLR(CLR), .D1(D[10]), .D2(D[11]), .EN1(EN), .EN2(EN),
           .PRE(gnd), .Q1(Q[10]), .Q2(Q[11]) );
dffepc_2 I5 ( .CLK(CLK), .CLR(CLR), .D1(D[8]), .D2(D[9]), .EN1(EN), .EN2(EN),
           .PRE(gnd), .Q1(Q[8]), .Q2(Q[9]) );
dffepc_2 I6 ( .CLK(CLK), .CLR(CLR), .D1(D[6]), .D2(D[7]), .EN1(EN), .EN2(EN),
           .PRE(gnd), .Q1(Q[6]), .Q2(Q[7]) );
dffepc_2 I7 ( .CLK(CLK), .CLR(CLR), .D1(D[4]), .D2(D[5]), .EN1(EN), .EN2(EN),
           .PRE(gnd), .Q1(Q[4]), .Q2(Q[5]) );
dffepc_2 I8 ( .CLK(CLK), .CLR(CLR), .D1(D[2]), .D2(D[3]), .EN1(EN), .EN2(EN),
           .PRE(gnd), .Q1(Q[2]), .Q2(Q[3]) );
dffepc_2 I9 ( .CLK(CLK), .CLR(CLR), .D1(D[0]), .D2(D[1]), .EN1(EN), .EN2(EN),
           .PRE(gnd), .Q1(Q[0]), .Q2(Q[1]) );

endmodule // rgec16_25um

`endif

`ifdef rge8_25um
`else
`define rge8_25um
module rge8_25um( CLK , D, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
 input [7:0] D;
input EN;
 output [7:0] Q;

dffe_2 I6 ( .CLK(CLK), .D1(D[6]), .D2(D[7]), .EN1(EN), .EN2(EN), .Q1(Q[6]),
         .Q2(Q[7]) );
dffe_2 I7 ( .CLK(CLK), .D1(D[4]), .D2(D[5]), .EN1(EN), .EN2(EN), .Q1(Q[4]),
         .Q2(Q[5]) );
dffe_2 I8 ( .CLK(CLK), .D1(D[2]), .D2(D[3]), .EN1(EN), .EN2(EN), .Q1(Q[2]),
         .Q2(Q[3]) );
dffe_2 I9 ( .CLK(CLK), .D1(D[0]), .D2(D[1]), .EN1(EN), .EN2(EN), .Q1(Q[0]),
         .Q2(Q[1]) );

endmodule // rge8_25um

`endif

`ifdef rge4_25um
`else
`define rge4_25um
module rge4_25um( CLK , D, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
 input [3:0] D;
input EN;
 output [3:0] Q;

dffe_2 I8 ( .CLK(CLK), .D1(D[2]), .D2(D[3]), .EN1(EN), .EN2(EN), .Q1(Q[2]),
         .Q2(Q[3]) );
dffe_2 I9 ( .CLK(CLK), .D1(D[0]), .D2(D[1]), .EN1(EN), .EN2(EN), .Q1(Q[0]),
         .Q2(Q[1]) );

endmodule // rge4_25um

`endif

`ifdef rge16_25um
`else
`define rge16_25um
module rge16_25um( CLK , D, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
 input [15:0] D;
input EN;
 output [15:0] Q;

dffe_2 I2 ( .CLK(CLK), .D1(D[14]), .D2(D[15]), .EN1(EN), .EN2(EN), .Q1(Q[14]),
         .Q2(Q[15]) );
dffe_2 I3 ( .CLK(CLK), .D1(D[12]), .D2(D[13]), .EN1(EN), .EN2(EN), .Q1(Q[12]),
         .Q2(Q[13]) );
dffe_2 I4 ( .CLK(CLK), .D1(D[10]), .D2(D[11]), .EN1(EN), .EN2(EN), .Q1(Q[10]),
         .Q2(Q[11]) );
dffe_2 I5 ( .CLK(CLK), .D1(D[8]), .D2(D[9]), .EN1(EN), .EN2(EN), .Q1(Q[8]),
         .Q2(Q[9]) );
dffe_2 I6 ( .CLK(CLK), .D1(D[6]), .D2(D[7]), .EN1(EN), .EN2(EN), .Q1(Q[6]),
         .Q2(Q[7]) );
dffe_2 I7 ( .CLK(CLK), .D1(D[4]), .D2(D[5]), .EN1(EN), .EN2(EN), .Q1(Q[4]),
         .Q2(Q[5]) );
dffe_2 I8 ( .CLK(CLK), .D1(D[2]), .D2(D[3]), .EN1(EN), .EN2(EN), .Q1(Q[2]),
         .Q2(Q[3]) );
dffe_2 I9 ( .CLK(CLK), .D1(D[0]), .D2(D[1]), .EN1(EN), .EN2(EN), .Q1(Q[0]),
         .Q2(Q[1]) );

endmodule // rge16_25um

`endif

`ifdef rgc8_25um
`else
`define rgc8_25um
module rgc8_25um( CLK , CLR, D, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [7:0] D;
 output [7:0] Q;

dffc_2 I6 ( .CLK(CLK), .CLR(CLR), .D1(D[6]), .D2(D[7]), .Q1(Q[6]), .Q2(Q[7]) );
dffc_2 I7 ( .CLK(CLK), .CLR(CLR), .D1(D[4]), .D2(D[5]), .Q1(Q[4]), .Q2(Q[5]) );
dffc_2 I8 ( .CLK(CLK), .CLR(CLR), .D1(D[0]), .D2(D[1]), .Q1(Q[0]), .Q2(Q[1]) );
dffc_2 I9 ( .CLK(CLK), .CLR(CLR), .D1(D[2]), .D2(D[3]), .Q1(Q[2]), .Q2(Q[3]) );

endmodule // rgc8_25um

`endif

`ifdef rgc4_25um
`else
`define rgc4_25um
module rgc4_25um( CLK , CLR, D, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [3:0] D;
 output [3:0] Q;

dffc_2 I8 ( .CLK(CLK), .CLR(CLR), .D1(D[0]), .D2(D[1]), .Q1(Q[0]), .Q2(Q[1]) );
dffc_2 I9 ( .CLK(CLK), .CLR(CLR), .D1(D[2]), .D2(D[3]), .Q1(Q[2]), .Q2(Q[3]) );

endmodule // rgc4_25um

`endif

`ifdef rgc16_25um
`else
`define rgc16_25um
module rgc16_25um( CLK , CLR, D, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [15:0] D;
 output [15:0] Q;

dffc_2 I2 ( .CLK(CLK), .CLR(CLR), .D1(D[14]), .D2(D[15]), .Q1(Q[14]), .Q2(Q[15]) );
dffc_2 I3 ( .CLK(CLK), .CLR(CLR), .D1(D[12]), .D2(D[13]), .Q1(Q[12]), .Q2(Q[13]) );
dffc_2 I4 ( .CLK(CLK), .CLR(CLR), .D1(D[10]), .D2(D[11]), .Q1(Q[10]), .Q2(Q[11]) );
dffc_2 I5 ( .CLK(CLK), .CLR(CLR), .D1(D[8]), .D2(D[9]), .Q1(Q[8]), .Q2(Q[9]) );
dffc_2 I6 ( .CLK(CLK), .CLR(CLR), .D1(D[6]), .D2(D[7]), .Q1(Q[6]), .Q2(Q[7]) );
dffc_2 I7 ( .CLK(CLK), .CLR(CLR), .D1(D[4]), .D2(D[5]), .Q1(Q[4]), .Q2(Q[5]) );
dffc_2 I8 ( .CLK(CLK), .CLR(CLR), .D1(D[0]), .D2(D[1]), .Q1(Q[0]), .Q2(Q[1]) );
dffc_2 I9 ( .CLK(CLK), .CLR(CLR), .D1(D[2]), .D2(D[3]), .Q1(Q[2]), .Q2(Q[3]) );

endmodule // rgc16_25um

`endif

`ifdef rg8_25um
`else
`define rg8_25um
module rg8_25um( CLK , D, Q );
input CLK /* synthesis syn_isclock=1 */;
 input [7:0] D;
 output [7:0] Q;

dff_2 I3 ( .CLK(CLK), .D1(D[6]), .D2(D[7]), .Q1(Q[6]), .Q2(Q[7]) );
dff_2 I4 ( .CLK(CLK), .D1(D[4]), .D2(D[5]), .Q1(Q[4]), .Q2(Q[5]) );
dff_2 I5 ( .CLK(CLK), .D1(D[0]), .D2(D[1]), .Q1(Q[0]), .Q2(Q[1]) );
dff_2 I6 ( .CLK(CLK), .D1(D[2]), .D2(D[3]), .Q1(Q[2]), .Q2(Q[3]) );

endmodule // rg8_25um

`endif

`ifdef rg4_25um
`else
`define rg4_25um
module rg4_25um( CLK , D, Q );
input CLK /* synthesis syn_isclock=1 */;
 input [3:0] D;
 output [3:0] Q;

dff_2 I3 ( .CLK(CLK), .D1(D[2]), .D2(D[3]), .Q1(Q[2]), .Q2(Q[3]) );
dff_2 I4 ( .CLK(CLK), .D1(D[0]), .D2(D[1]), .Q1(Q[0]), .Q2(Q[1]) );

endmodule // rg4_25um

`endif

`ifdef rg16_25um
`else
`define rg16_25um
module rg16_25um( CLK , D, Q );
input CLK /* synthesis syn_isclock=1 */;
 input [15:0] D;
 output [15:0] Q;

dff_2 I6 ( .CLK(CLK), .D1(D[14]), .D2(D[15]), .Q1(Q[14]), .Q2(Q[15]) );
dff_2 I7 ( .CLK(CLK), .D1(D[12]), .D2(D[13]), .Q1(Q[12]), .Q2(Q[13]) );
dff_2 I8 ( .CLK(CLK), .D1(D[10]), .D2(D[11]), .Q1(Q[10]), .Q2(Q[11]) );
dff_2 I9 ( .CLK(CLK), .D1(D[8]), .D2(D[9]), .Q1(Q[8]), .Q2(Q[9]) );
dff_2 I2 ( .CLK(CLK), .D1(D[6]), .D2(D[7]), .Q1(Q[6]), .Q2(Q[7]) );
dff_2 I3 ( .CLK(CLK), .D1(D[4]), .D2(D[5]), .Q1(Q[4]), .Q2(Q[5]) );
dff_2 I4 ( .CLK(CLK), .D1(D[2]), .D2(D[3]), .Q1(Q[2]), .Q2(Q[3]) );
dff_2 I5 ( .CLK(CLK), .D1(D[0]), .D2(D[1]), .Q1(Q[0]), .Q2(Q[1]) );

endmodule // rg16_25um

`endif

`ifdef dffepc_2
`else
`define dffepc_2
module dffepc_2( CLK , CLR, D1, D2, EN1, EN2, PRE, Q1, Q2 );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input PRE /* synthesis syn_isclock=1 */;
input D1, D2, EN1, EN2;
output Q1, Q2;
supply1 vcc;
supply0 gnd;

super_logic I4 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(gnd),
              .B1(Q1), .B2(gnd), .C1(D1), .C2(gnd), .D1(Q2), .D2(gnd), .E1(D2),
              .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd), .F5(vcc),
              .F6(gnd), .MP(gnd), .MS(EN1), .NP(gnd), .NS(EN2), .OP(gnd),
              .OS(gnd), .PP(gnd), .PS(gnd), .Q2Z(Q2), .QC(CLK), .QR(CLR),
              .QS(PRE), .QZ(Q1) );

endmodule // dffepc_2

`endif

`ifdef dffe_2
`else
`define dffe_2
module dffe_2( CLK , D1, D2, EN1, EN2, Q1, Q2 );
input CLK /* synthesis syn_isclock=1 */;
input D1, D2, EN1, EN2;
output Q1, Q2;
supply0 gnd;
supply1 vcc;

super_logic I2 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(gnd),
              .B1(Q1), .B2(gnd), .C1(D1), .C2(gnd), .D1(Q2), .D2(gnd), .E1(D2),
              .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd), .F5(vcc),
              .F6(gnd), .MP(gnd), .MS(EN1), .NP(gnd), .NS(EN2), .OP(gnd),
              .OS(gnd), .PP(gnd), .PS(gnd), .Q2Z(Q2), .QC(CLK), .QR(gnd),
              .QS(gnd), .QZ(Q1) );

endmodule // dffe_2

`endif

`ifdef dffc_2
`else
`define dffc_2
module dffc_2( CLK , CLR, D1, D2, Q1, Q2 );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input D1, D2;
output Q1, Q2;
supply1 vcc;
supply0 gnd;

super_logic I3 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(gnd),
              .B1(vcc), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd),
              .E1(D1), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd),
              .F5(vcc), .F6(gnd), .MP(gnd), .MS(gnd), .NP(gnd), .NS(vcc),
              .OP(gnd), .OS(vcc), .PP(vcc), .PS(D2), .Q2Z(Q2), .QC(CLK),
              .QR(CLR), .QS(gnd), .QZ(Q1) );

endmodule // dffc_2

`endif

`ifdef dff_2
`else
`define dff_2
module dff_2( CLK , D1, D2, Q1, Q2 );
input CLK /* synthesis syn_isclock=1 */;
input D1, D2;
output Q1, Q2;
supply1 vcc;
supply0 gnd;

super_logic I2 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(gnd),
              .B1(vcc), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd),
              .E1(D1), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd),
              .F5(vcc), .F6(gnd), .MP(gnd), .MS(vcc), .NP(gnd), .NS(vcc),
              .OP(gnd), .OS(vcc), .PP(vcc), .PS(D2), .Q2Z(Q2), .QC(CLK),
              .QR(gnd), .QS(gnd), .QZ(Q1) );

endmodule // dff_2

`endif

`ifdef super_logic
`else
`define super_logic
module super_logic( A1 , A2, A3, A4, A5, A6, B1, B2, C1, C2, D1, D2, E1, E2, F1,
                    F2, F3, F4, F5, F6, MP, MS, NP, NS, OP, OS, PP, PS, QC,
                    QR, QS, AZ, FZ, NZ, OZ, Q2Z, QZ );
input A1, A2, A3, A4, A5, A6;
output AZ;
input B1, B2, C1, C2, D1, D2, E1, E2, F1, F2, F3, F4, F5, F6;
output FZ;
input MP, MS, NP, NS;
output NZ;
input OP, OS;
output OZ;
input PP, PS;
output Q2Z;
input QC /* synthesis syn_isclock=1 */;
input QR /* synthesis syn_isclock=1 */;
input QS /* synthesis syn_isclock=1 */;
output QZ;
parameter ql_gate = `LOGIC;

super_cell I2 ( .A1(A1), .A2(A2), .A3(A3), .A4(A4), .A5(A5), .A6(A6), .AZ(AZ),
             .B1(B1), .B2(B2), .C1(C1), .C2(C2), .D1(D1), .D2(D2), .E1(E1),
             .E2(E2), .F1(F1), .F2(F2), .F3(F3), .F4(F4), .F5(F5), .F6(F6),
             .FZ(FZ), .MP(MP), .MS(MS), .NP(NP), .NS(NS), .NZ(NZ), .OP(OP),
             .OS(OS), .OZ(OZ), .PP(PP), .PS(PS), .Q2Z(Q2Z), .QC(QC), .QR(QR),
             .QS(QS), .QZ(QZ) );

endmodule // super_logic

`endif

`ifdef gclkbuff_25um
`else
`define gclkbuff_25um
module gclkbuff_25um( A , Z );
input A;
output Z;
parameter ql_gate = `HSCKMUX;
supply1 vcc;

hsckmux I1 ( .IC(A), .IS(vcc), .IZ(Z) );

endmodule // gclkbuff_25um

`endif

`ifdef inv_gclkbuff_25um
`else
`define inv_gclkbuff_25um
module inv_gclkbuff_25um( A , Z );
input A;
output Z;
supply1 vcc;
supply0 gnd;
wire N_1;

super_logic I1 ( .A1(vcc), .A2(A), .A3(vcc), .A4(gnd), .A5(vcc), .A6(gnd), .AZ(N_1),
              .B1(gnd), .B2(gnd), .C1(gnd), .C2(gnd), .D1(gnd), .D2(gnd),
              .E1(gnd), .E2(gnd), .F1(gnd), .F2(gnd), .F3(gnd), .F4(gnd),
              .F5(gnd), .F6(gnd), .MP(gnd), .MS(gnd), .NP(gnd), .NS(gnd),
              .OP(gnd), .OS(gnd), .PP(gnd), .PS(gnd), .QC(gnd), .QR(gnd),
              .QS(vcc) );
gclkbuff_25um I2 ( .A(N_1), .Z(Z) );

endmodule // inv_gclkbuff_25um

`endif


`ifdef tripados_25um
`else
`define tripados_25um
module tripados_25um( EN , P );
input EN;
output P;
parameter ql_gate = `BIDIR;
supply0 GND;
supply1 VCC;

eio_cell I1 ( .EQE(VCC), .ESEL(VCC), .IE(EN), .IP(P), .IQC(GND), .IQE(GND),
           .IQR(GND), .OQI(VCC), .OSEL(VCC) );

endmodule // tripados_25um

`endif

`ifdef tripadod_25um
`else
`define tripadod_25um
module tripadod_25um( EN , P );
input EN;
output P;
parameter ql_gate = `BIDIR;
supply0 GND;
supply1 VCC;

eio_cell I3 ( .EQE(VCC), .ESEL(VCC), .IE(EN), .IP(P), .IQC(GND), .IQE(GND),
           .IQR(GND), .OQI(GND), .OSEL(VCC) );

endmodule // tripadod_25um

`endif

`ifdef tripadff_25um
`else
`define tripadff_25um
module tripadff_25um( A , EN, FFCLK, FFCLR, P, Q );
input A, EN;
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
output P, Q;
parameter ql_gate = `BIDIR;
supply0 GND;
supply1 VCC;

eio_cell I1 ( .EQE(VCC), .ESEL(VCC), .IE(EN), .IP(P), .IQC(FFCLK), .IQE(GND),
           .IQR(FFCLR), .IZ(Q), .OQI(A), .OSEL(GND) );

endmodule // tripadff_25um

`endif

`ifdef tripad_25um
`else
`define tripad_25um
module tripad_25um( A , EN, P );
input A, EN;
output P;
parameter ql_gate = `BIDIR;
supply0 GND;
supply1 VCC;

eio_cell I1 ( .EQE(VCC), .ESEL(VCC), .IE(EN), .IP(P), .IQC(GND), .IQE(GND),
           .IQR(GND), .OQI(A), .OSEL(VCC) );

endmodule // tripad_25um

`endif

`ifdef outpadff_25um
`else
`define outpadff_25um
module outpadff_25um( A , FFCLK, FFCLR, P, P_FB );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input A;
output P, P_FB;
parameter ql_gate = `BIDIR;
supply0 GND;
supply1 VCC;

eio_cell I1 ( .EQE(VCC), .ESEL(VCC), .IE(VCC), .IP(P), .IQC(FFCLK), .IQE(GND),
           .IQR(FFCLR), .OQI(A), .OQQ(P_FB), .OSEL(GND) );

endmodule // outpadff_25um

`endif

`ifdef outpad_25um
`else
`define outpad_25um
module outpad_25um( A , P );
input A;
output P;
parameter ql_gate = `BIDIR;
supply0 GND;
supply1 VCC;

eio_cell I1 ( .EQE(VCC), .ESEL(VCC), .IE(VCC), .IP(P), .IQC(GND), .IQE(GND),
           .IQR(GND), .OQI(A), .OSEL(VCC) );

endmodule // outpad_25um

`endif

`ifdef inpadff_25um
`else
`define inpadff_25um
module inpadff_25um( FFCLK , FFCLR, FFEN, P, FFQ, Q );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input FFEN;
output FFQ;
input P;
output Q;
parameter ql_gate = `BIDIR;
supply0 gnd;
supply1 vcc;

eio_cell I1 ( .EQE(vcc), .ESEL(vcc), .IE(gnd), .IP(P), .IQC(FFCLK), .IQE(FFEN),
           .IQQ(FFQ), .IQR(FFCLR), .IZ(Q), .OQI(gnd), .OSEL(vcc) );

endmodule // inpadff_25um

`endif

`ifdef io_buff_25um
`else
`define io_buff_25um
module io_buff_25um( I , O );
input I;
output O;
parameter ql_gate = `IOCONTROL;
supply0 gnd;
supply1 vcc;

inbuffcell_25um I1 ( .I(I), .IP(gnd), .IS(vcc), .O(O) );

endmodule // io_buff_25um

`endif

`ifdef inpad_25um
`else
`define inpad_25um
module inpad_25um( P , Q );
input P;
output Q;
parameter ql_gate = `BIDIR;
supply0 gnd;
supply1 vcc;

eio_cell I1 ( .EQE(vcc), .ESEL(vcc), .IE(gnd), .IP(P), .IQC(gnd), .IQE(gnd),
           .IQR(gnd), .IZ(Q), .OQI(vcc), .OSEL(vcc) );

endmodule // inpad_25um

`endif

`ifdef hdpad_25um
`else
`define hdpad_25um
module hdpad_25um( IP , O );
input IP;
output O;
parameter ql_gate = `IOCONTROL;
supply0 gnd;

iocontrol I1 ( .IP(IP), .IS(GND), .O(O) );

endmodule // hdpad_25um

`endif

`ifdef eio_25um
`else
`define eio_25um
module eio_25um( A2 , EN, FFCLK, FFCLR, I_EN, OE_EN, OESEL, OSEL, FFQ, P_FB, Q,
                 P );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input A2, EN;
output FFQ;
input I_EN, OE_EN, OESEL, OSEL;
inout P;
output P_FB, Q;
parameter ql_gate = `BIDIR;

eio_cell I1 ( .EQE(OE_EN), .ESEL(OESEL), .IE(EN), .IP(P), .IQC(FFCLK), .IQE(I_EN),
           .IQQ(FFQ), .IQR(FFCLR), .IZ(Q), .OQI(A2), .OQQ(P_FB), .OSEL(OSEL) );

endmodule // eio_25um

`endif

`ifdef ckpad_25um
`else
`define ckpad_25um
module ckpad_25um( P , Q );
input P /*synthesis syn_isclock=1 */;
output Q;
parameter ql_gate = `CLOCK;

ckcell_25um I1 ( .IC(Q), .IP(P) );

endmodule // ckpad_25um

`endif

`ifdef bipados_25um
`else
`define bipados_25um
module bipados_25um( EN , Q, P );
input EN;
inout P;
output Q;
parameter ql_gate = `BIDIR;
supply0 gnd;
supply1 vcc;

eio_cell I1 ( .EQE(vcc), .ESEL(vcc), .IE(EN), .IP(P), .IQC(gnd), .IQE(gnd),
           .IQR(gnd), .IZ(Q), .OQI(vcc), .OSEL(vcc) );

endmodule // bipados_25um

`endif

`ifdef bipadoff_25um
`else
`define bipadoff_25um
module bipadoff_25um( A2 , EN, FFCLK, FFCLR, P_FB, Q, P );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input A2, EN;
inout P;
output P_FB, Q;
parameter ql_gate = `BIDIR;
supply0 gnd;
supply1 vcc;

eio_cell I1 ( .EQE(vcc), .ESEL(vcc), .IE(EN), .IP(P), .IQC(FFCLK), .IQE(gnd),
           .IQR(FFCLR), .IZ(Q), .OQI(A2), .OQQ(P_FB), .OSEL(gnd) );

endmodule // bipadoff_25um

`endif

`ifdef bipadod_25um
`else
`define bipadod_25um
module bipadod_25um( EN , Q, P );
input EN;
inout P;
output Q;
parameter ql_gate = `BIDIR;
supply0 gnd;
supply1 vcc;

eio_cell I1 ( .EQE(vcc), .ESEL(vcc), .IE(EN), .IP(P), .IQC(gnd), .IQE(gnd),
           .IQR(gnd), .IZ(Q), .OQI(gnd), .OSEL(vcc) );

endmodule // bipadod_25um

`endif

`ifdef bipadioff_25um
`else
`define bipadioff_25um
module bipadioff_25um( A2 , EN, FFCLK, FFCLR, inFFEN, FFQ, P_FB, Q, P );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input A2, EN;
output FFQ;
input inFFEN;
inout P;
output P_FB, Q;
parameter ql_gate = `BIDIR;
supply0 gnd;
supply1 vcc;

eio_cell I1 ( .EQE(vcc), .ESEL(vcc), .IE(EN), .IP(P), .IQC(FFCLK), .IQE(inFFEN),
           .IQQ(FFQ), .IQR(FFCLR), .IZ(Q), .OQI(A2), .OQQ(P_FB), .OSEL(gnd) );

endmodule // bipadioff_25um

`endif

`ifdef bipadiff_25um
`else
`define bipadiff_25um
module bipadiff_25um( A2 , EN, FFCLK, FFCLR, FFEN, FFQ, Q, P );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input FFEN;
input A2, EN;
output FFQ;
inout P;
output Q;
parameter ql_gate = `BIDIR;
supply1 vcc;

eio_cell I1 ( .EQE(vcc), .ESEL(vcc), .IE(EN), .IP(P), .IQC(FFCLK), .IQE(FFEN),
           .IQQ(FFQ), .IQR(FFCLR), .IZ(Q), .OQI(A2), .OSEL(vcc) );

endmodule // bipadiff_25um

`endif

`ifdef bipadeioff_25um
`else
`define bipadeioff_25um
module bipadeioff_25um( A2 , EN, FFCLK, FFCLR, I_EN, OE_EN, FFQ, P_FB, Q, P );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input A2, EN;
output FFQ;
input I_EN, OE_EN;
inout P;
output P_FB, Q;
parameter ql_gate = `BIDIR;
supply0 gnd;

eio_cell I1 ( .EQE(OE_EN), .ESEL(gnd), .IE(EN), .IP(P), .IQC(FFCLK), .IQE(I_EN),
           .IQQ(FFQ), .IQR(FFCLR), .IZ(Q), .OQI(A2), .OQQ(P_FB), .OSEL(gnd) );

endmodule // bipadeioff_25um

`endif

`ifdef bipad_25um
`else
`define bipad_25um
module bipad_25um( A , EN, Q, P );
input A, EN;
inout P;
output Q;
parameter ql_gate = `BIDIR;
supply0 gnd;
supply1 vcc;

eio_cell I2 ( .EQE(vcc), .ESEL(vcc), .IE(EN), .IP(P), .IQC(gnd), .IQE(gnd),
           .IQR(gnd), .IZ(Q), .OQI(A), .OSEL(vcc) );

endmodule // bipad_25um

`endif

`ifdef ckpadp5
`else
`define ckpadp5
module ckpadp5( P , Q );
input P /*synthesis syn_isclock=1 */;
output Q;
parameter ql_gate = `CLOCKB;

ckcell5 I3 ( .IC(Q), .IP(P) );

endmodule // ckpadp5

`endif

`ifdef ucebitb0
`else
`define ucebitb0
module ucebitb0( CLK , CLR, ENH1, ENH2, ENH3, ENH4, ENL1, ENL2, ENL3, QFB, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input ENH1, ENH2, ENH3, ENH4, ENL1, ENL2, ENL3;
output Q;
input QFB;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

lcell2 I_1 ( .A1(ENH2), .A2(ENL3), .A3(ENH3), .A4(ENL2), .A5(ENH4), .A6(ENL1),
          .B1(GND), .B2(GND), .C1(VCC), .C2(QFB), .D1(QFB), .D2(GND), .E1(GND),
          .E2(GND), .F1(VCC), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND),
          .MP(GND), .MS(VCC), .NP(GND), .NS(GND), .OP(ENH1), .OS(GND), .QC(CLK),
          .QR(CLR), .QS(GND), .QZ(Q) );

endmodule // ucebitb0

`endif

`ifdef udrn6_p2
`else
`define udrn6_p2
module udrn6_p2( ARST , CLK, D, D0, D1, D2N, DOWN, LDN, Q, U0, U1, U2N, UPN,
                 ALLONEN, ALLZERO );
output ALLONEN, ALLZERO;
input CLK /* synthesis syn_isclock=1 */;
input ARST;
 input [5:0] D;
input D0, D1, D2N, DOWN, LDN;
 input [5:0] Q;
input U0, U1, U2N, UPN;
wire N_15;
wire N_16;
wire N_12;
wire N_14;
wire N_9;
wire N_10;
wire N_7;
supply1 VCC;
supply0 GND;

or2i0 I_12 ( .A(ALLONEN), .B(N_16), .Q(N_15) );
and5i3 I_10 ( .A(U0), .B(U1), .C(DOWN), .D(U2N), .E(UPN), .Q(N_12) );
and5i2 I_11 ( .A(DOWN), .B(UPN), .C(D2N), .D(D1), .E(D0), .Q(N_16) );
and16i7 I_5 ( .A(VCC), .B(VCC), .C(VCC), .D(VCC), .E(VCC), .F(VCC), .G(D2N), .H(UPN),
           .I(DOWN), .J(D1), .K(D0), .L(Q[1]), .M(Q[2]), .N(Q[3]), .O(Q[4]),
           .P(Q[5]), .Q(N_7) );
and16i7 I_6 ( .A(Q[1]), .B(Q[2]), .C(Q[3]), .D(Q[4]), .E(Q[5]), .F(U0), .G(U1),
           .H(VCC), .I(VCC), .J(UPN), .K(DOWN), .L(U2N), .M(GND), .N(GND),
           .O(GND), .P(GND), .Q(N_14) );
logic2 I_8 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .B1(VCC),
          .B2(VCC), .C1(GND), .C2(GND), .D1(GND), .D2(VCC), .E1(D[5]), .E2(GND),
          .F1(D[3]), .F2(GND), .F3(D[2]), .F4(GND), .F5(D[1]), .F6(GND),
          .MP(GND), .MS(GND), .NP(D[4]), .NS(GND), .OP(GND), .OS(D[0]), .OZ(N_9),
          .QC(GND), .QR(GND), .QS(GND) );
logic2 I_3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(D[0]), .A5(VCC), .A6(D[5]), .B1(GND),
          .B2(GND), .C1(VCC), .C2(VCC), .D1(VCC), .D2(VCC), .E1(VCC), .E2(D[4]),
          .F1(VCC), .F2(D[3]), .F3(VCC), .F4(D[2]), .F5(VCC), .F6(D[1]),
          .MP(GND), .MS(GND), .NP(VCC), .NS(GND), .OP(VCC), .OS(GND), .OZ(N_10),
          .QC(GND), .QR(GND), .QS(GND) );
logic2 I_7 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .B1(VCC),
          .B2(N_9), .C1(VCC), .C2(VCC), .D1(Q[0]), .D2(GND), .E1(N_15), .E2(GND),
          .F1(VCC), .F2(N_14), .F3(VCC), .F4(N_7), .F5(VCC), .F6(GND), .MP(GND),
          .MS(GND), .NP(VCC), .NS(GND), .OP(GND), .OS(LDN), .QC(CLK), .QR(GND),
          .QS(ARST), .QZ(ALLONEN) );
logic2 I_1 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .B1(N_10),
          .B2(GND), .C1(VCC), .C2(VCC), .D1(Q[0]), .D2(GND), .E1(ALLZERO),
          .E2(N_12), .F1(VCC), .F2(N_14), .F3(VCC), .F4(N_7), .F5(VCC), .F6(GND),
          .MP(GND), .MS(GND), .NP(VCC), .NS(GND), .OP(GND), .OS(LDN), .QC(CLK),
          .QR(GND), .QS(ARST), .QZ(ALLZERO) );

endmodule // udrn6_p2

`endif

`ifdef udrc6_p2
`else
`define udrc6_p2
module udrc6_p2( ARST , CLK, D, D0, D1, D2N, DOWN, LDN, Q, U0, U1, U2N, UPN,
                 ALLONE, ALLZERON );
output ALLONE, ALLZERON;
input CLK /* synthesis syn_isclock=1 */;
input ARST;
 input [5:0] D;
input D0, D1, D2N, DOWN, LDN;
 input [5:0] Q;
input U0, U1, U2N, UPN;
wire N_13;
wire N_14;
wire N_12;
wire N_7;
wire N_8;
wire N_6;
supply1 VCC;
supply0 GND;
wire N_1;

or2i0 I_13 ( .A(N_14), .B(ALLZERON), .Q(N_13) );
and5i2 I_12 ( .A(DOWN), .B(UPN), .C(D2N), .D(D1), .E(D0), .Q(N_12) );
and5i3 I_11 ( .A(U0), .B(U1), .C(DOWN), .D(U2N), .E(UPN), .Q(N_14) );
and16i7 I_6 ( .A(Q[1]), .B(Q[2]), .C(Q[3]), .D(Q[4]), .E(Q[5]), .F(U0), .G(U1),
           .H(VCC), .I(VCC), .J(UPN), .K(DOWN), .L(U2N), .M(GND), .N(GND),
           .O(GND), .P(GND), .Q(N_8) );
and16i7 I_5 ( .A(VCC), .B(VCC), .C(VCC), .D(VCC), .E(VCC), .F(VCC), .G(D2N), .H(UPN),
           .I(DOWN), .J(D1), .K(D0), .L(Q[1]), .M(Q[2]), .N(Q[3]), .O(Q[4]),
           .P(Q[5]), .Q(N_7) );
logic2 I_7 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .B1(N_6),
          .B2(GND), .C1(VCC), .C2(VCC), .D1(VCC), .D2(Q[0]), .E1(ALLONE),
          .E2(N_12), .F1(VCC), .F2(N_8), .F3(VCC), .F4(N_7), .F5(VCC), .F6(GND),
          .MP(GND), .MS(GND), .NP(VCC), .NS(GND), .OP(GND), .OS(LDN), .QC(CLK),
          .QR(ARST), .QS(GND), .QZ(ALLONE) );
logic2 I_8 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .B1(VCC),
          .B2(VCC), .C1(GND), .C2(GND), .D1(GND), .D2(VCC), .E1(D[5]), .E2(GND),
          .F1(D[3]), .F2(GND), .F3(D[2]), .F4(GND), .F5(D[1]), .F6(GND),
          .MP(GND), .MS(GND), .NP(D[4]), .NS(GND), .OP(GND), .OS(D[0]), .OZ(N_6),
          .QC(GND), .QR(GND), .QS(GND) );
logic2 I_1 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .B1(VCC),
          .B2(N_1), .C1(VCC), .C2(VCC), .D1(VCC), .D2(Q[0]), .E1(N_13), .E2(GND),
          .F1(VCC), .F2(N_8), .F3(VCC), .F4(N_7), .F5(VCC), .F6(GND), .MP(GND),
          .MS(GND), .NP(VCC), .NS(GND), .OP(GND), .OS(LDN), .QC(CLK), .QR(ARST),
          .QS(GND), .QZ(ALLZERON) );
logic2 I_3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(D[0]), .A5(VCC), .A6(D[5]), .B1(GND),
          .B2(GND), .C1(VCC), .C2(VCC), .D1(VCC), .D2(VCC), .E1(VCC), .E2(D[4]),
          .F1(VCC), .F2(D[3]), .F3(VCC), .F4(D[2]), .F5(VCC), .F6(D[1]),
          .MP(GND), .MS(GND), .NP(VCC), .NS(GND), .OP(VCC), .OS(GND), .OZ(N_1),
          .QC(GND), .QR(GND), .QS(GND) );

endmodule // udrc6_p2

`endif

`ifdef udlf6
`else
`define udlf6
module udlf6( ARST , CLK, D, DOWN, LDN, UPN, MAX, MIN, Q );
input CLK /* synthesis syn_isclock=1 */;
input ARST;
 input [5:0] D;
input DOWN, LDN;
output MAX, MIN;
 output [5:0] Q;
input UPN;
wire RCDN1;
supply0 GND;
supply1 VCC;

inv I_24 ( .A(RCDN1), .Q(MIN) );
ud6fs_p2 I_21 ( .ARST(ARST), .CLK(CLK), .D({ D[5:0] }), .D0(GND), .D1(GND),
             .D3N(VCC), .DOWN(DOWN), .LDN(LDN), .Q({ Q[5:0] }), .U0(VCC),
             .U1(VCC), .U3N(GND), .UPN(UPN) );
udrc6_p2 I_17 ( .ALLONE(MAX), .ALLZERON(RCDN1), .ARST(ARST), .CLK(CLK),
             .D({ D[5:0] }), .D0(GND), .D1(GND), .D2N(VCC), .DOWN(DOWN),
             .LDN(LDN), .Q({ Q[5:0] }), .U0(VCC), .U1(VCC), .U2N(GND),
             .UPN(UPN) );

endmodule // udlf6

`endif

`ifdef udlf24
`else
`define udlf24
module udlf24( ARST , CLK, D, DOWN, LDN, UPN, MAX, MIN, Q );
input CLK /* synthesis syn_isclock=1 */;
input ARST;
 input [23:0] D;
input DOWN, LDN;
output MAX, MIN;
 output [23:0] Q;
input UPN;
wire LDNB;
wire RCUN4;
wire RCUN3;
wire RCD4;
wire RCD3;
supply0 GND;
supply1 VCC;
wire RCDN2;
wire RCU2;
wire RCDN1;
wire RCU1;

ud6fs_p2 I_18 ( .ARST(ARST), .CLK(CLK), .D({ D[23:18] }), .D0(RCDN1), .D1(RCDN2),
             .D3N(RCD3), .DOWN(DOWN), .LDN(LDN), .Q({ Q[23:18] }), .U0(RCU1),
             .U1(RCU2), .U3N(RCUN3), .UPN(UPN) );
ud6fs_p2 I_19 ( .ARST(ARST), .CLK(CLK), .D({ D[17:12] }), .D0(RCDN1), .D1(RCDN2),
             .D3N(VCC), .DOWN(DOWN), .LDN(LDN), .Q({ Q[17:12] }), .U0(RCU1),
             .U1(RCU2), .U3N(GND), .UPN(UPN) );
ud6fs_p2 I_20 ( .ARST(ARST), .CLK(CLK), .D({ D[11:6] }), .D0(RCDN1), .D1(GND),
             .D3N(VCC), .DOWN(DOWN), .LDN(LDN), .Q({ Q[11:6] }), .U0(RCU1),
             .U1(VCC), .U3N(GND), .UPN(UPN) );
ud6fs_p2 I_21 ( .ARST(ARST), .CLK(CLK), .D({ D[5:0] }), .D0(GND), .D1(GND),
             .D3N(VCC), .DOWN(DOWN), .LDN(LDN), .Q({ Q[5:0] }), .U0(VCC),
             .U1(VCC), .U3N(GND), .UPN(UPN) );
and4i2 I_12 ( .A(RCD4), .B(RCD3), .C(RCDN2), .D(RCDN1), .Q(MIN) );
and4i2 I_13 ( .A(RCU1), .B(RCU2), .C(RCUN3), .D(RCUN4), .Q(MAX) );
udrn6_p2 I_15 ( .ALLONEN(RCUN3), .ALLZERO(RCD3), .ARST(ARST), .CLK(CLK),
             .D({ D[17:12] }), .D0(RCDN1), .D1(RCDN2), .D2N(VCC), .DOWN(DOWN),
             .LDN(LDNB), .Q({ Q[17:12] }), .U0(RCU1), .U1(RCU2), .U2N(GND),
             .UPN(UPN) );
udrn6_p2 I_14 ( .ALLONEN(RCUN4), .ALLZERO(RCD4), .ARST(ARST), .CLK(CLK),
             .D({ D[23:18] }), .D0(RCDN1), .D1(RCDN2), .D2N(RCD3), .DOWN(DOWN),
             .LDN(LDNB), .Q({ Q[23:18] }), .U0(RCU1), .U1(RCU2), .U2N(RCUN3),
             .UPN(UPN) );
udrc6_p2 I_17 ( .ALLONE(RCU1), .ALLZERON(RCDN1), .ARST(ARST), .CLK(CLK),
             .D({ D[5:0] }), .D0(GND), .D1(GND), .D2N(VCC), .DOWN(DOWN),
             .LDN(LDNB), .Q({ Q[5:0] }), .U0(VCC), .U1(VCC), .U2N(GND),
             .UPN(UPN) );
udrc6_p2 I_16 ( .ALLONE(RCU2), .ALLZERON(RCDN2), .ARST(ARST), .CLK(CLK),
             .D({ D[11:6] }), .D0(RCDN1), .D1(GND), .D2N(VCC), .DOWN(DOWN),
             .LDN(LDNB), .Q({ Q[11:6] }), .U0(RCU1), .U1(VCC), .U2N(GND),
             .UPN(UPN) );
buff I_11 ( .A(LDN), .Q(LDNB) );

endmodule // udlf24

`endif

`ifdef udlf18
`else
`define udlf18
module udlf18( ARST , CLK, D, DOWN, LDN, UPN, MAX, MIN, Q );
input CLK /* synthesis syn_isclock=1 */;
input ARST;
 input [17:0] D;
input DOWN, LDN;
output MAX, MIN;
 output [17:0] Q;
input UPN;
wire LDNB;
wire RCUN3;
wire RCD3;
supply0 GND;
supply1 VCC;
wire RCDN2;
wire RCU2;
wire RCDN1;
wire RCU1;

and3i2 I_22 ( .A(RCD3), .B(RCDN2), .C(RCDN1), .Q(MIN) );
and3i1 I_23 ( .A(RCU1), .B(RCU2), .C(RCUN3), .Q(MAX) );
ud6fs_p2 I_19 ( .ARST(ARST), .CLK(CLK), .D({ D[17:12] }), .D0(RCDN1), .D1(RCDN2),
             .D3N(VCC), .DOWN(DOWN), .LDN(LDN), .Q({ Q[17:12] }), .U0(RCU1),
             .U1(RCU2), .U3N(GND), .UPN(UPN) );
ud6fs_p2 I_20 ( .ARST(ARST), .CLK(CLK), .D({ D[11:6] }), .D0(RCDN1), .D1(GND),
             .D3N(VCC), .DOWN(DOWN), .LDN(LDN), .Q({ Q[11:6] }), .U0(RCU1),
             .U1(VCC), .U3N(GND), .UPN(UPN) );
ud6fs_p2 I_21 ( .ARST(ARST), .CLK(CLK), .D({ D[5:0] }), .D0(GND), .D1(GND),
             .D3N(VCC), .DOWN(DOWN), .LDN(LDN), .Q({ Q[5:0] }), .U0(VCC),
             .U1(VCC), .U3N(GND), .UPN(UPN) );
udrn6_p2 I_15 ( .ALLONEN(RCUN3), .ALLZERO(RCD3), .ARST(ARST), .CLK(CLK),
             .D({ D[17:12] }), .D0(RCDN1), .D1(RCDN2), .D2N(VCC), .DOWN(DOWN),
             .LDN(LDNB), .Q({ Q[17:12] }), .U0(RCU1), .U1(RCU2), .U2N(GND),
             .UPN(UPN) );
udrc6_p2 I_17 ( .ALLONE(RCU1), .ALLZERON(RCDN1), .ARST(ARST), .CLK(CLK),
             .D({ D[5:0] }), .D0(GND), .D1(GND), .D2N(VCC), .DOWN(DOWN),
             .LDN(LDNB), .Q({ Q[5:0] }), .U0(VCC), .U1(VCC), .U2N(GND),
             .UPN(UPN) );
udrc6_p2 I_16 ( .ALLONE(RCU2), .ALLZERON(RCDN2), .ARST(ARST), .CLK(CLK),
             .D({ D[11:6] }), .D0(RCDN1), .D1(GND), .D2N(VCC), .DOWN(DOWN),
             .LDN(LDNB), .Q({ Q[11:6] }), .U0(RCU1), .U1(VCC), .U2N(GND),
             .UPN(UPN) );
buff I_11 ( .A(LDN), .Q(LDNB) );

endmodule // udlf18

`endif

`ifdef udlf12
`else
`define udlf12
module udlf12( ARST , CLK, D, DOWN, LDN, UPN, MAX, MIN, Q );
input CLK /* synthesis syn_isclock=1 */;
input ARST;
 input [11:0] D;
input DOWN, LDN;
output MAX, MIN;
 output [11:0] Q;
input UPN;
wire LDNB;
supply0 GND;
supply1 VCC;
wire RCDN2;
wire RCU2;
wire RCDN1;
wire RCU1;

and2i2 I_23 ( .A(RCDN1), .B(RCDN2), .Q(MIN) );
and2i0 I_24 ( .A(RCU1), .B(RCU2), .Q(MAX) );
ud6fs_p2 I_20 ( .ARST(ARST), .CLK(CLK), .D({ D[11:6] }), .D0(RCDN1), .D1(GND),
             .D3N(VCC), .DOWN(DOWN), .LDN(LDN), .Q({ Q[11:6] }), .U0(RCU1),
             .U1(VCC), .U3N(GND), .UPN(UPN) );
ud6fs_p2 I_21 ( .ARST(ARST), .CLK(CLK), .D({ D[5:0] }), .D0(GND), .D1(GND),
             .D3N(VCC), .DOWN(DOWN), .LDN(LDN), .Q({ Q[5:0] }), .U0(VCC),
             .U1(VCC), .U3N(GND), .UPN(UPN) );
udrc6_p2 I_17 ( .ALLONE(RCU1), .ALLZERON(RCDN1), .ARST(ARST), .CLK(CLK),
             .D({ D[5:0] }), .D0(GND), .D1(GND), .D2N(VCC), .DOWN(DOWN),
             .LDN(LDNB), .Q({ Q[5:0] }), .U0(VCC), .U1(VCC), .U2N(GND),
             .UPN(UPN) );
udrc6_p2 I_16 ( .ALLONE(RCU2), .ALLZERON(RCDN2), .ARST(ARST), .CLK(CLK),
             .D({ D[11:6] }), .D0(RCDN1), .D1(GND), .D2N(VCC), .DOWN(DOWN),
             .LDN(LDNB), .Q({ Q[11:6] }), .U0(RCU1), .U1(VCC), .U2N(GND),
             .UPN(UPN) );
buff I_11 ( .A(LDN), .Q(LDNB) );

endmodule // udlf12

`endif

`ifdef udbtb_p2
`else
`define udbtb_p2
module udbtb_p2( ARST , CLK, D, D0, D1, D2, D3N, D4N, D5N, LDN, U0, U1, U2, U3N,
                 U4N, U5N, DE, Q, UE );
input CLK /* synthesis syn_isclock=1 */;
input ARST, D, D0, D1, D2, D3N, D4N, D5N;
output DE;
input LDN;
output Q;
input U0, U1, U2, U3N, U4N, U5N;
output UE;
parameter syn_macro = 1, ql_pack = 1;
supply1 VCC;
supply0 GND;

logic2 I_1 ( .A1(U0), .A2(U3N), .A3(U1), .A4(U4N), .A5(U2), .A6(U5N), .AZ(UE),
          .B1(Q), .B2(GND), .C1(VCC), .C2(Q), .D1(VCC), .D2(Q), .E1(D), .E2(GND),
          .F1(D5N), .F2(D0), .F3(D4N), .F4(D1), .F5(D3N), .F6(D2), .FZ(DE),
          .MP(VCC), .MS(GND), .NP(LDN), .NS(VCC), .OP(LDN), .OS(VCC), .QC(CLK),
          .QR(ARST), .QS(GND), .QZ(Q) );

endmodule // udbtb_p2

`endif

`ifdef ud6fs_p2
`else
`define ud6fs_p2
module ud6fs_p2( ARST , CLK, D, D0, D1, D3N, DOWN, LDN, U0, U1, U3N, UPN, Q );
input CLK /* synthesis syn_isclock=1 */;
input ARST;
 input [5:0] D;
input D0, D1, D3N, DOWN, LDN;
 output [5:0] Q;
input U0, U1, U3N, UPN;
wire LDNB;
supply1 VCC;
wire UE0;
wire Q2N;
wire Q1N;
wire Q0N;
wire DE0;
supply0 GND;

buff I_11 ( .A(LDN), .Q(LDNB) );
inv I_8 ( .A(Q[2]), .Q(Q2N) );
inv I_9 ( .A(Q[1]), .Q(Q1N) );
inv I_10 ( .A(Q[0]), .Q(Q0N) );
udbtb_p2 BIT5 ( .ARST(ARST), .CLK(CLK), .D(D[5]), .D0(Q[0]), .D1(Q[4]), .D2(Q[3]),
             .D3N(Q2N), .D4N(Q1N), .D5N(DE0), .LDN(LDNB), .Q(Q[5]), .U0(UE0),
             .U1(Q[4]), .U2(Q[3]), .U3N(Q2N), .U4N(Q1N), .U5N(Q0N) );
udbtb_p2 BIT4 ( .ARST(ARST), .CLK(CLK), .D(D[4]), .D0(Q[1]), .D1(Q[3]), .D2(GND),
             .D3N(Q2N), .D4N(DE0), .D5N(Q0N), .LDN(LDNB), .Q(Q[4]), .U0(UE0),
             .U1(Q[3]), .U2(VCC), .U3N(Q2N), .U4N(Q1N), .U5N(Q0N) );
udbtb_p2 BIT3 ( .ARST(ARST), .CLK(CLK), .D(D[3]), .D0(Q[2]), .D1(GND), .D2(GND),
             .D3N(DE0), .D4N(Q1N), .D5N(Q0N), .LDN(LDNB), .Q(Q[3]), .U0(UE0),
             .U1(VCC), .U2(VCC), .U3N(Q2N), .U4N(Q1N), .U5N(Q0N) );
udbtb_p2 BIT2 ( .ARST(ARST), .CLK(CLK), .D(D[2]), .D0(GND), .D1(GND), .D2(GND),
             .D3N(Q1N), .D4N(Q0N), .D5N(DE0), .LDN(LDNB), .Q(Q[2]), .U0(UE0),
             .U1(VCC), .U2(VCC), .U3N(Q1N), .U4N(Q0N), .U5N(GND) );
udbtb_p2 BIT1 ( .ARST(ARST), .CLK(CLK), .D(D[1]), .D0(GND), .D1(GND), .D2(GND),
             .D3N(Q0N), .D4N(VCC), .D5N(DE0), .LDN(LDNB), .Q(Q[1]), .U0(UE0),
             .U1(VCC), .U2(VCC), .U3N(Q0N), .U4N(GND), .U5N(GND) );
udbtb_p2 BIT0 ( .ARST(ARST), .CLK(CLK), .D(D[0]), .D0(D0), .D1(D1), .D2(GND),
             .D3N(D3N), .D4N(UPN), .D5N(DOWN), .DE(DE0), .LDN(LDNB), .Q(Q[0]),
             .U0(U0), .U1(U1), .U2(VCC), .U3N(U3N), .U4N(DOWN), .U5N(UPN),
             .UE(UE0) );

endmodule // ud6fs_p2

`endif

`ifdef uctx16p2
`else
`define uctx16p2
module uctx16p2( CLK , CLR, D, EN, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [15:0] D;
input EN, LOAD;
 output [15:0] Q;
wire UCTXCO;
wire Q8BUFFN1;
wire Q3Q4Q5EN1;
wire Q3EN;
wire Q13BUFFN1;
wire Q12BUFFN1;
wire Q4BUFF1;
wire Q0BUFF1;
wire D0D1D2;
wire Q1Q2Q0N;
wire LDBUFFN3;
wire Q3Q4Q5EN2;
wire Q6Q7Q8;
wire Q9Q10Q11;
wire Q7BUFFN1;
wire Q6BUFF1;
wire LDBUFFN2;
wire ENBUFF1;
wire LDBUFFN1;
wire CO3;
wire CO2;
supply1 VCC;
supply0 GND;
wire CO1;

ucxco UCXCO1 ( .CLK(CLK), .CO(UCTXCO), .D_DEC(D0D1D2), .EN(ENBUFF1),
            .LDBUF(LDBUFFN1), .LOAD(LOAD), .PRE(CLR), .Q_DEC(Q1Q2Q0N) );
and4i1 I_90 ( .A(Q[3]), .B(Q[4]), .C(Q[5]), .D(EN), .Q(Q3Q4Q5EN1) );
and4i1 I_94 ( .A(Q[7]), .B(Q[6]), .C(Q[8]), .D(EN), .Q(Q3Q4Q5EN2) );
ucxbit2b UCTX8 ( .CLK(CLK), .CLR(CLR), .D(D[8]), .ENH1(Q3Q4Q5EN1), .ENH2(Q6BUFF1),
              .ENH3(VCC), .ENH4(VCC), .ENL1(CO2), .ENL2(Q7BUFFN1), .ENL3(GND),
              .LOAD(LDBUFFN2), .Q(Q[8]), .QFB(Q8BUFFN1) );
ucxbit2b UCTX13 ( .CLK(CLK), .CLR(CLR), .D(D[13]), .ENH1(Q3Q4Q5EN2),
               .ENH2(Q6Q7Q8), .ENH3(Q9Q10Q11), .ENH4(VCC), .ENL1(CO3),
               .ENL2(Q12BUFFN1), .ENL3(GND), .LOAD(LDBUFFN3), .Q(Q[13]),
               .QFB(Q13BUFFN1) );
ucxbit2b UCTX12 ( .CLK(CLK), .CLR(CLR), .D(D[12]), .ENH1(Q3Q4Q5EN2),
               .ENH2(Q6Q7Q8), .ENH3(Q9Q10Q11), .ENH4(VCC), .ENL1(CO3),
               .ENL2(GND), .ENL3(GND), .LOAD(LDBUFFN3), .Q(Q[12]),
               .QFB(Q12BUFFN1) );
ucxbit2b UCTX7 ( .CLK(CLK), .CLR(CLR), .D(D[7]), .ENH1(Q3EN), .ENH2(Q4BUFF1),
              .ENH3(Q[5]), .ENH4(Q6BUFF1), .ENL1(CO1), .ENL2(GND), .ENL3(GND),
              .LOAD(LDBUFFN2), .Q(Q[7]), .QFB(Q7BUFFN1) );
ucxbit2a UCTX14 ( .CLK(CLK), .CLR(CLR), .D(D[14]), .ENH1(Q3Q4Q5EN2),
               .ENH2(Q6Q7Q8), .ENH3(Q9Q10Q11), .ENH4(VCC), .ENL1(CO3),
               .ENL2(Q12BUFFN1), .ENL3(Q13BUFFN1), .LOAD(LDBUFFN3), .Q(Q[14]),
               .QFB(Q[14]) );
ucxbit2a UCTX15 ( .CLK(CLK), .CLR(CLR), .D(D[15]), .ENH1(Q3Q4Q5EN2),
               .ENH2(Q6Q7Q8), .ENH3(Q9Q10Q11), .ENH4(Q[14]), .ENL1(CO3),
               .ENL2(Q12BUFFN1), .ENL3(Q13BUFFN1), .LOAD(LDBUFFN3), .Q(Q[15]),
               .QFB(Q[15]) );
ucxbit2a UCTX4 ( .CLK(CLK), .CLR(CLR), .D(D[4]), .ENH1(Q3EN), .ENH2(VCC),
              .ENH3(VCC), .ENH4(VCC), .ENL1(CO1), .ENL2(GND), .ENL3(GND),
              .LOAD(LDBUFFN2), .Q(Q[4]), .QFB(Q4BUFF1) );
ucxbit2a UCTX5 ( .CLK(CLK), .CLR(CLR), .D(D[5]), .ENH1(Q3EN), .ENH2(Q4BUFF1),
              .ENH3(VCC), .ENH4(VCC), .ENL1(CO1), .ENL2(GND), .ENL3(GND),
              .LOAD(LDBUFFN2), .Q(Q[5]), .QFB(Q[5]) );
ucxbit2a UCTX9 ( .CLK(CLK), .CLR(CLR), .D(D[9]), .ENH1(Q3Q4Q5EN1), .ENH2(Q6BUFF1),
              .ENH3(VCC), .ENH4(VCC), .ENL1(CO2), .ENL2(Q7BUFFN1),
              .ENL3(Q8BUFFN1), .LOAD(LDBUFFN2), .Q(Q[9]), .QFB(Q[9]) );
ucxbit2a UCTX10 ( .CLK(CLK), .CLR(CLR), .D(D[10]), .ENH1(Q3Q4Q5EN1),
               .ENH2(Q6BUFF1), .ENH3(Q[9]), .ENH4(VCC), .ENL1(CO2),
               .ENL2(Q7BUFFN1), .ENL3(Q8BUFFN1), .LOAD(LDBUFFN3), .Q(Q[10]),
               .QFB(Q[10]) );
ucxbit2a UCTX6 ( .CLK(CLK), .CLR(CLR), .D(D[6]), .ENH1(Q3EN), .ENH2(Q4BUFF1),
              .ENH3(Q[5]), .ENH4(VCC), .ENL1(CO1), .ENL2(GND), .ENL3(GND),
              .LOAD(LDBUFFN2), .Q(Q[6]), .QFB(Q6BUFF1) );
ucxbit2a UCTX11 ( .CLK(CLK), .CLR(CLR), .D(D[11]), .ENH1(Q3Q4Q5EN1),
               .ENH2(Q6BUFF1), .ENH3(Q[9]), .ENH4(Q[10]), .ENL1(CO2),
               .ENL2(Q7BUFFN1), .ENL3(Q8BUFFN1), .LOAD(LDBUFFN3), .Q(Q[11]),
               .QFB(Q[11]) );
ucxbit2a UCTX3 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENH1(Q0BUFF1), .ENH2(Q[1]),
              .ENH3(Q[2]), .ENH4(VCC), .ENL1(ENBUFF1), .ENL2(GND), .ENL3(GND),
              .LOAD(LDBUFFN1), .Q(Q[3]), .QFB(Q[3]) );
ucxbit2a UCTX2 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENH1(Q0BUFF1), .ENH2(Q[1]),
              .ENH3(VCC), .ENH4(VCC), .ENL1(ENBUFF1), .ENL2(GND), .ENL3(GND),
              .LOAD(LDBUFFN1), .Q(Q[2]), .QFB(Q[2]) );
ucxbit2a UCTX1 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENH1(Q0BUFF1), .ENH2(VCC),
              .ENH3(VCC), .ENH4(VCC), .ENL1(ENBUFF1), .ENL2(GND), .ENL3(GND),
              .LOAD(LDBUFFN1), .Q(Q[1]), .QFB(Q[1]) );
ucxbit2a UCTX0 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENH1(VCC), .ENH2(VCC),
              .ENH3(VCC), .ENH4(VCC), .ENL1(ENBUFF1), .ENL2(GND), .ENL3(GND),
              .LOAD(LDBUFFN1), .Q(Q[0]), .QFB(Q0BUFF1) );
and3i0 I_95 ( .A(Q[9]), .B(Q[10]), .C(Q[11]), .Q(Q9Q10Q11) );
and3i0 I_96 ( .A(Q[3]), .B(Q[4]), .C(Q[5]), .Q(Q6Q7Q8) );
and3i0 I_104 ( .A(D[0]), .B(D[1]), .C(D[2]), .Q(D0D1D2) );
inv I_34 ( .A(Q[7]), .Q(Q7BUFFN1) );
inv I_99 ( .A(Q[13]), .Q(Q13BUFFN1) );
inv I_100 ( .A(Q[12]), .Q(Q12BUFFN1) );
inv I_92 ( .A(Q[8]), .Q(Q8BUFFN1) );
inv I_111 ( .A(LOAD), .Q(LDBUFFN3) );
inv I_107 ( .A(LOAD), .Q(LDBUFFN2) );
and3i1 I_105 ( .A(Q[1]), .B(Q[2]), .C(Q[0]), .Q(Q1Q2Q0N) );
and2i1 I_72 ( .A(Q[3]), .B(EN), .Q(Q3EN) );
buff I_93 ( .A(Q[6]), .Q(Q6BUFF1) );
buff I_42 ( .A(Q[4]), .Q(Q4BUFF1) );
buff I_32 ( .A(Q[0]), .Q(Q0BUFF1) );
buff I_112 ( .A(UCTXCO), .Q(CO1) );
buff I_114 ( .A(UCTXCO), .Q(CO3) );
buff I_113 ( .A(UCTXCO), .Q(CO2) );
buff I_108 ( .A(EN), .Q(ENBUFF1) );

endmodule // uctx16p2

`endif

`ifdef ucte16p2
`else
`define ucte16p2
module ucte16p2( CLK , CLR, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input EN;
 output [15:0] Q;
wire Q1Q2Q3;
wire UCTECO;
wire Q11BUFFN1;
wire Q10Q13;
wire Q12BUFFN1;
wire Q7Q8Q9;
wire Q4Q5Q6EN1;
wire Q4Q5Q6EN2;
wire Q8BUFFN1;
wire Q10BUFF1;
wire Q7BUFF1;
wire ENBUFFN2;
wire Q5BUFF1;
wire Q4BUFF1;
wire Q0BUFF1;
supply0 GND;
wire ENBUFFN1;
wire CO1A;
supply1 VCC;
wire CO1B;
wire CO1C;
wire N_13;

and2i0 I_62 ( .A(Q[10]), .B(Q[13]), .Q(Q10Q13) );
ucebit2b UCTE12 ( .CLK(CLK), .CLR(CLR), .ENH1(Q4Q5Q6EN2), .ENH2(Q7Q8Q9),
               .ENH3(Q10BUFF1), .ENH4(VCC), .ENL1(CO1C), .ENL2(GND),
               .ENL3(Q11BUFFN1), .Q(Q[12]), .QFB(Q12BUFFN1) );
ucebit2b UCTE8 ( .CLK(CLK), .CLR(CLR), .ENH1(Q4Q5Q6EN1), .ENH2(Q7BUFF1),
              .ENH3(VCC), .ENH4(VCC), .ENL1(CO1B), .ENL2(GND), .ENL3(GND),
              .Q(Q[8]), .QFB(Q8BUFFN1) );
mux4x2 I_34 ( .A(VCC), .B(Q[0]), .C(VCC), .D(Q[0]), .Q(N_13), .S0(Q1Q2Q3),
           .S1(ENBUFFN1) );
inv I_44 ( .A(Q[11]), .Q(Q11BUFFN1) );
inv I_58 ( .A(Q[12]), .Q(Q12BUFFN1) );
inv I_57 ( .A(Q[8]), .Q(Q8BUFFN1) );
inv I_56 ( .A(EN), .Q(ENBUFFN2) );
inv I_35 ( .A(EN), .Q(ENBUFFN1) );
and4i1 I_45 ( .A(Q[4]), .B(Q[5]), .C(Q[6]), .D(EN), .Q(Q4Q5Q6EN2) );
and4i1 I_59 ( .A(Q[4]), .B(Q[5]), .C(Q[6]), .D(EN), .Q(Q4Q5Q6EN1) );
buff I_33 ( .A(UCTECO), .Q(CO1A) );
buff I_47 ( .A(UCTECO), .Q(CO1C) );
buff I_32 ( .A(UCTECO), .Q(CO1B) );
buff I_60 ( .A(Q[7]), .Q(Q7BUFF1) );
buff I_63 ( .A(Q[10]), .Q(Q10BUFF1) );
buff I_51 ( .A(Q[4]), .Q(Q4BUFF1) );
buff I_50 ( .A(Q[5]), .Q(Q5BUFF1) );
buff I_49 ( .A(Q[0]), .Q(Q0BUFF1) );
and3i0 I_17 ( .A(Q[1]), .B(Q[2]), .C(Q[3]), .Q(Q1Q2Q3) );
and3i0 I_61 ( .A(Q[7]), .B(Q[8]), .C(Q[9]), .Q(Q7Q8Q9) );
dffp I_18 ( .CLK(CLK), .D(N_13), .PRE(CLR), .Q(UCTECO) );
ucebit2a UCTE15 ( .CLK(CLK), .CLR(CLR), .ENH1(Q4Q5Q6EN2), .ENH2(Q7Q8Q9),
               .ENH3(Q10Q13), .ENH4(Q[14]), .ENL1(CO1C), .ENL2(Q11BUFFN1),
               .ENL3(Q12BUFFN1), .Q(Q[15]), .QFB(Q[15]) );
ucebit2a UCTE14 ( .CLK(CLK), .CLR(CLR), .ENH1(Q4Q5Q6EN2), .ENH2(Q7Q8Q9),
               .ENH3(Q10Q13), .ENH4(VCC), .ENL1(CO1C), .ENL2(Q11BUFFN1),
               .ENL3(Q12BUFFN1), .Q(Q[14]), .QFB(Q[14]) );
ucebit2a UCTE13 ( .CLK(CLK), .CLR(CLR), .ENH1(Q4Q5Q6EN2), .ENH2(Q7Q8Q9),
               .ENH3(Q10BUFF1), .ENH4(VCC), .ENL1(CO1C), .ENL2(Q11BUFFN1),
               .ENL3(Q12BUFFN1), .Q(Q[13]), .QFB(Q[13]) );
ucebit2a UCTE11 ( .CLK(CLK), .CLR(CLR), .ENH1(Q4Q5Q6EN1), .ENH2(Q7BUFF1),
               .ENH3(Q[9]), .ENH4(Q10BUFF1), .ENL1(CO1B), .ENL2(Q8BUFFN1),
               .ENL3(GND), .Q(Q[11]), .QFB(Q[11]) );
ucebit2a UCTE10 ( .CLK(CLK), .CLR(CLR), .ENH1(Q4Q5Q6EN1), .ENH2(Q7BUFF1),
               .ENH3(Q[9]), .ENH4(VCC), .ENL1(CO1B), .ENL2(Q8BUFFN1),
               .ENL3(GND), .Q(Q[10]), .QFB(Q10BUFF1) );
ucebit2a UCTE9 ( .CLK(CLK), .CLR(CLR), .ENH1(Q4Q5Q6EN1), .ENH2(Q7BUFF1),
              .ENH3(VCC), .ENH4(VCC), .ENL1(CO1B), .ENL2(Q8BUFFN1), .ENL3(GND),
              .Q(Q[9]), .QFB(Q[9]) );
ucebit2a UCTE7 ( .CLK(CLK), .CLR(CLR), .ENH1(ENBUFFN2), .ENH2(Q4BUFF1),
              .ENH3(Q5BUFF1), .ENH4(Q[6]), .ENL1(CO1A), .ENL2(GND), .ENL3(GND),
              .Q(Q[7]), .QFB(Q[7]) );
ucebit2a UCTE6 ( .CLK(CLK), .CLR(CLR), .ENH1(ENBUFFN2), .ENH2(Q4BUFF1),
              .ENH3(Q5BUFF1), .ENH4(VCC), .ENL1(CO1A), .ENL2(GND), .ENL3(GND),
              .Q(Q[6]), .QFB(Q[6]) );
ucebit2a UCTE5 ( .CLK(CLK), .CLR(CLR), .ENH1(ENBUFFN2), .ENH2(Q4BUFF1),
              .ENH3(VCC), .ENH4(VCC), .ENL1(CO1A), .ENL2(GND), .ENL3(GND),
              .Q(Q[5]), .QFB(Q5BUFF1) );
ucebit2a UCTE4 ( .CLK(CLK), .CLR(CLR), .ENH1(ENBUFFN2), .ENH2(VCC), .ENH3(VCC),
              .ENH4(VCC), .ENL1(CO1A), .ENL2(GND), .ENL3(GND), .Q(Q[4]),
              .QFB(Q4BUFF1) );
ucebit2a UCTE3 ( .CLK(CLK), .CLR(CLR), .ENH1(ENBUFFN1), .ENH2(Q0BUFF1),
              .ENH3(Q[1]), .ENH4(Q[2]), .ENL1(GND), .ENL2(GND), .ENL3(GND),
              .Q(Q[3]), .QFB(Q[3]) );
ucebit2a UCTE2 ( .CLK(CLK), .CLR(CLR), .ENH1(ENBUFFN1), .ENH2(Q0BUFF1),
              .ENH3(Q[1]), .ENH4(VCC), .ENL1(GND), .ENL2(GND), .ENL3(GND),
              .Q(Q[2]), .QFB(Q[2]) );
ucebit2a UCTE1 ( .CLK(CLK), .CLR(CLR), .ENH1(ENBUFFN1), .ENH2(Q0BUFF1),
              .ENH3(VCC), .ENH4(VCC), .ENL1(GND), .ENL2(GND), .ENL3(GND),
              .Q(Q[1]), .QFB(Q[1]) );
ucebit2a UCTE0 ( .CLK(CLK), .CLR(CLR), .ENH1(ENBUFFN1), .ENH2(VCC), .ENH3(VCC),
              .ENH4(VCC), .ENL1(GND), .ENL2(GND), .ENL3(GND), .Q(Q[0]),
              .QFB(Q0BUFF1) );

endmodule // ucte16p2

`endif

`ifdef sub32p2
`else
`define sub32p2
module sub32p2( A , B, Bi, Bo, Diff );
 input [31:0] A;
 input [31:0] B;
input Bi;
output Bo;
 output [31:0] Diff;
wire [31:0] S;
wire Carry15;
wire Carry15a;
wire Carry15b;
wire Co0_Ci0;
wire Co0_Ci1;
wire Co1_C00;
wire Co1_C01;
wire Co2_C10;
wire Co2_C11;
wire Co3_C20;
wire Co3_C21;
wire Co4_C30;
wire Co4_C31;
wire Co5_C40;
wire Co5_C41;
wire Co6_C50;
wire Co6_C51;
wire Co8_C70;
wire Co8_C71;
wire Co9_C80;
wire Co9_C81;
wire Co10_C90;
wire Co10_C91;
wire Co12_C110;
wire Co12_C111;
wire Co13_C120;
wire Co13_C121;
wire Co14_C130;
wire Co14_C131;
wire Co16_C150;
wire Co16_C151;
wire Co17_C160;
wire Carry3;
wire Co17_C161;
wire Carry3a;
wire Co18_C170;
wire Co18_C171;
wire Co20_C190;
wire Co20_C191;
wire Co21_C200;
wire Co21_C201;
wire Co22_C210;
wire Co22_C211;
wire Co24_C230;
wire Co24_C231;
wire Co25_C240;
wire Co25_C241;
wire Co26_C250;
wire Co26_C251;
wire Co28_C270;
wire Co28_C271;
wire Co29_C280;
wire Co29_C281;
wire Co30_C290;
wire Co30_C291;
wire C7_C30;
wire C7_C31;
wire C11_C70;
wire C11_C71;
wire C19_C150;
wire C19_C151;
wire C23_C190;
wire C23_C191;
wire C27_C230;
wire C27_C231;

dif32 I_7 ( .a({ A[0] }), .b({ B[0] }), .C11_C70(C11_C70), .C11_C71(C11_C71),
         .C19_C150(C19_C150), .C19_C151(C19_C151), .C23_C190(C23_C190),
         .C23_C191(C23_C191), .C27_C230(C27_C230), .C27_C231(C27_C231),
         .C7_C30(C7_C30), .C7_C31(C7_C31), .Carry15(Carry15),
         .Carry15a(Carry15a), .Carry15b(Carry15b), .Carry3(Carry3),
         .Carry3a(Carry3a), .Cin(Bi), .Co0_Ci0(Co0_Ci0), .Co0_Ci1(Co0_Ci1),
         .Co10_C90(Co10_C90), .Co10_C91(Co10_C91), .Co12_C110(Co12_C110),
         .Co12_C111(Co12_C111), .Co13_C120(Co13_C120), .Co13_C121(Co13_C121),
         .Co14_C130(Co14_C130), .Co14_C131(Co14_C131), .Co16_C150(Co16_C150),
         .Co16_C151(Co16_C151), .Co17_C160(Co17_C160), .Co17_C161(Co17_C161),
         .Co18_C170(Co18_C170), .Co18_C171(Co18_C171), .Co1_C00(Co1_C00),
         .Co1_C01(Co1_C01), .Co20_C190(Co20_C190), .Co20_C191(Co20_C191),
         .Co21_C200(Co21_C200), .Co21_C201(Co21_C201), .Co22_C210(Co22_C210),
         .Co22_C211(Co22_C211), .Co24_C230(Co24_C230), .Co24_C231(Co24_C231),
         .Co25_C240(Co25_C240), .Co25_C241(Co25_C241), .Co26_C250(Co26_C250),
         .Co26_C251(Co26_C251), .Co28_C270(Co28_C270), .Co28_C271(Co28_C271),
         .Co29_C280(Co29_C280), .Co29_C281(Co29_C281), .Co2_C10(Co2_C10),
         .Co2_C11(Co2_C11), .Co30_C290(Co30_C290), .Co30_C291(Co30_C291),
         .Co3_C20(Co3_C20), .Co3_C21(Co3_C21), .Co4_C30(Co4_C30),
         .Co4_C31(Co4_C31), .Co5_C40(Co5_C40), .Co5_C41(Co5_C41),
         .Co6_C50(Co6_C50), .Co6_C51(Co6_C51), .Co8_C70(Co8_C70),
         .Co8_C71(Co8_C71), .Co9_C80(Co9_C80), .Co9_C81(Co9_C81),
         .S({ S[31:0] }), .Sumi({ Diff[31:0] }) );
borrow32 I_6 ( .a({ A[31:0] }), .b({ B[31:0] }), .C11_C70(C11_C70),
            .C11_C71(C11_C71), .C19_C150(C19_C150), .C19_C151(C19_C151),
            .C23_C190(C23_C190), .C23_C191(C23_C191), .C27_C230(C27_C230),
            .C27_C231(C27_C231), .C7_C30(C7_C30), .C7_C31(C7_C31),
            .Carry15(Carry15), .Carry15a(Carry15a), .Carry15b(Carry15b),
            .Carry3(Carry3), .Carry3a(Carry3a), .Co(Bo), .Co0_Ci0(Co0_Ci0),
            .Co0_Ci1(Co0_Ci1), .Co10_C90(Co10_C90), .Co10_C91(Co10_C91),
            .Co12_C110(Co12_C110), .Co12_C111(Co12_C111),
            .Co13_C120(Co13_C120), .Co13_C121(Co13_C121),
            .Co14_C130(Co14_C130), .Co14_C131(Co14_C131),
            .Co16_C150(Co16_C150), .Co16_C151(Co16_C151),
            .Co17_C160(Co17_C160), .Co17_C161(Co17_C161),
            .Co18_C170(Co18_C170), .Co18_C171(Co18_C171), .Co1_C00(Co1_C00),
            .Co1_C01(Co1_C01), .Co20_C190(Co20_C190), .Co20_C191(Co20_C191),
            .Co21_C200(Co21_C200), .Co21_C201(Co21_C201),
            .Co22_C210(Co22_C210), .Co22_C211(Co22_C211),
            .Co24_C230(Co24_C230), .Co24_C231(Co24_C231),
            .Co25_C240(Co25_C240), .Co25_C241(Co25_C241),
            .Co26_C250(Co26_C250), .Co26_C251(Co26_C251),
            .Co28_C270(Co28_C270), .Co28_C271(Co28_C271),
            .Co29_C280(Co29_C280), .Co29_C281(Co29_C281), .Co2_C10(Co2_C10),
            .Co2_C11(Co2_C11), .Co30_C290(Co30_C290), .Co30_C291(Co30_C291),
            .Co3_C20(Co3_C20), .Co3_C21(Co3_C21), .Co4_C30(Co4_C30),
            .Co4_C31(Co4_C31), .Co5_C40(Co5_C40), .Co5_C41(Co5_C41),
            .Co6_C50(Co6_C50), .Co6_C51(Co6_C51), .Co8_C70(Co8_C70),
            .Co8_C71(Co8_C71), .Co9_C80(Co9_C80), .Co9_C81(Co9_C81),
            .S({ S[31:0] }) );

endmodule // sub32p2

`endif

`ifdef sub16p2
`else
`define sub16p2
module sub16p2( A , B, Bi, Bo, Diff );
 input [15:0] A;
 input [15:0] B;
input Bi;
output Bo;
 output [15:0] Diff;
wire [15:0] D;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire Borrow3;
wire Co0_Ci0;
wire Co0_Ci1;
wire Co1_C00;
wire Co1_C01;
wire Co2_C10;
wire Co2_C11;
wire Co3_C20;
wire Co3_C21;
wire Co4_C30;
wire Co4_C31;
wire Co5_C40;
wire Co5_C41;
wire Co6_C50;
wire Co6_C51;
wire Co8_C70;
wire Co8_C71;
wire Co9_C80;
wire Co9_C81;
wire Co10_C90;
wire Co10_C91;
wire Co12_C110;
wire Co12_C111;
wire Co13_C120;
wire Co13_C121;
wire Co14_C130;
wire Co14_C131;

borrow16 I_10 ( .a({ A[15:0] }), .b({ B[15:0] }), .Bo(Bo), .Borrow3(Borrow3),
             .C11_C70(N_3), .C11_C71(N_2), .C7_C30(N_5), .C7_C31(N_4),
             .Co0_Ci0(Co0_Ci0), .Co0_Ci1(Co0_Ci1), .Co10_C90(Co10_C90),
             .Co10_C91(Co10_C91), .Co12_C110(Co12_C110),
             .Co12_C111(Co12_C111), .Co13_C120(Co13_C120),
             .Co13_C121(Co13_C121), .Co14_C130(Co14_C130),
             .Co14_C131(Co14_C131), .Co1_C00(Co1_C00), .Co1_C01(Co1_C01),
             .Co2_C10(Co2_C10), .Co2_C11(Co2_C11), .Co3_C20(Co3_C20),
             .Co3_C21(Co3_C21), .Co4_C30(Co4_C30), .Co4_C31(Co4_C31),
             .Co5_C40(Co5_C40), .Co5_C41(Co5_C41), .Co6_C50(Co6_C50),
             .Co6_C51(Co6_C51), .Co8_C70(Co8_C70), .Co8_C71(Co8_C71),
             .Co9_C80(Co9_C80), .Co9_C81(Co9_C81), .D({ D[15:0] }) );
dif16 I_9 ( .a({ A[0] }), .b({ B[0] }), .Bin(Bi), .Borrow3(Borrow3),
         .C11_C70(N_3), .C11_C71(N_2), .C7_C30(N_5), .C7_C31(N_4),
         .Co0_Ci0(Co0_Ci0), .Co0_Ci1(Co0_Ci1), .Co10_C90(Co10_C90),
         .Co10_C91(Co10_C91), .Co12_C110(Co12_C110), .Co12_C111(Co12_C111),
         .Co13_C120(Co13_C120), .Co13_C121(Co13_C121), .Co14_C130(Co14_C130),
         .Co14_C131(Co14_C131), .Co1_C00(Co1_C00), .Co1_C01(Co1_C01),
         .Co2_C10(Co2_C10), .Co2_C11(Co2_C11), .Co3_C20(Co3_C20),
         .Co3_C21(Co3_C21), .Co4_C30(Co4_C30), .Co4_C31(Co4_C31),
         .Co5_C40(Co5_C40), .Co5_C41(Co5_C41), .Co6_C50(Co6_C50),
         .Co6_C51(Co6_C51), .Co8_C70(Co8_C70), .Co8_C71(Co8_C71),
         .Co9_C80(Co9_C80), .Co9_C81(Co9_C81), .D({ D[15:0] }),
         .Diffi({ Diff[15:0] }) );

endmodule // sub16p2

`endif

`ifdef add32p2
`else
`define add32p2
module add32p2( A , B, Ci, Co, Sum );
 input [31:0] A;
 input [31:0] B;
input Ci;
output Co;
 output [31:0] Sum;
wire [31:0] S;
wire Carry15;
wire Carry15a;
wire Carry15b;
wire Co0_Ci0;
wire Co0_Ci1;
wire Co1_C00;
wire Co1_C01;
wire Co2_C10;
wire Co2_C11;
wire Co3_C20;
wire Co3_C21;
wire Co4_C30;
wire Co4_C31;
wire Co5_C40;
wire Co5_C41;
wire Co6_C50;
wire Co6_C51;
wire Co8_C70;
wire Co8_C71;
wire Co9_C80;
wire Co9_C81;
wire Co10_C90;
wire Co10_C91;
wire Co12_C110;
wire Co12_C111;
wire Co13_C120;
wire Co13_C121;
wire Co14_C130;
wire Co14_C131;
wire Co16_C150;
wire Co16_C151;
wire Co17_C160;
wire Carry3;
wire Co17_C161;
wire Carry3a;
wire Co18_C170;
wire Co18_C171;
wire Co20_C190;
wire Co20_C191;
wire Co21_C200;
wire Co21_C201;
wire Co22_C210;
wire Co22_C211;
wire Co24_C230;
wire Co24_C231;
wire Co25_C240;
wire Co25_C241;
wire Co26_C250;
wire Co26_C251;
wire Co28_C270;
wire Co28_C271;
wire Co29_C280;
wire Co29_C281;
wire Co30_C290;
wire Co30_C291;
wire C7_C30;
wire C7_C31;
wire C11_C70;
wire C11_C71;
wire C19_C150;
wire C19_C151;
wire C23_C190;
wire C23_C191;
wire C27_C230;
wire C27_C231;

carry32 I2 ( .a({ A[31:0] }), .b({ B[31:0] }), .C11_C70(C11_C70),
          .C11_C71(C11_C71), .C19_C150(C19_C150), .C19_C151(C19_C151),
          .C23_C190(C23_C190), .C23_C191(C23_C191), .C27_C230(C27_C230),
          .C27_C231(C27_C231), .C7_C30(C7_C30), .C7_C31(C7_C31),
          .Carry15(Carry15), .Carry15a(Carry15a), .Carry15b(Carry15b),
          .Carry3(Carry3), .Carry3a(Carry3a), .Co(Co), .Co0_Ci0(Co0_Ci0),
          .Co0_Ci1(Co0_Ci1), .Co10_C90(Co10_C90), .Co10_C91(Co10_C91),
          .Co12_C110(Co12_C110), .Co12_C111(Co12_C111),
          .Co13_C120(Co13_C120), .Co13_C121(Co13_C121),
          .Co14_C130(Co14_C130), .Co14_C131(Co14_C131),
          .Co16_C150(Co16_C150), .Co16_C151(Co16_C151),
          .Co17_C160(Co17_C160), .Co17_C161(Co17_C161),
          .Co18_C170(Co18_C170), .Co18_C171(Co18_C171), .Co1_C00(Co1_C00),
          .Co1_C01(Co1_C01), .Co20_C190(Co20_C190), .Co20_C191(Co20_C191),
          .Co21_C200(Co21_C200), .Co21_C201(Co21_C201),
          .Co22_C210(Co22_C210), .Co22_C211(Co22_C211),
          .Co24_C230(Co24_C230), .Co24_C231(Co24_C231),
          .Co25_C240(Co25_C240), .Co25_C241(Co25_C241),
          .Co26_C250(Co26_C250), .Co26_C251(Co26_C251),
          .Co28_C270(Co28_C270), .Co28_C271(Co28_C271),
          .Co29_C280(Co29_C280), .Co29_C281(Co29_C281), .Co2_C10(Co2_C10),
          .Co2_C11(Co2_C11), .Co30_C290(Co30_C290), .Co30_C291(Co30_C291),
          .Co3_C20(Co3_C20), .Co3_C21(Co3_C21), .Co4_C30(Co4_C30),
          .Co4_C31(Co4_C31), .Co5_C40(Co5_C40), .Co5_C41(Co5_C41),
          .Co6_C50(Co6_C50), .Co6_C51(Co6_C51), .Co8_C70(Co8_C70),
          .Co8_C71(Co8_C71), .Co9_C80(Co9_C80), .Co9_C81(Co9_C81),
          .S({ S[31:0] }) );
sum32 I3 ( .a({ A[0] }), .b({ B[0] }), .C11_C70(C11_C70), .C11_C71(C11_C71),
        .C19_C150(C19_C150), .C19_C151(C19_C151), .C23_C190(C23_C190),
        .C23_C191(C23_C191), .C27_C230(C27_C230), .C27_C231(C27_C231),
        .C7_C30(C7_C30), .C7_C31(C7_C31), .Carry15(Carry15),
        .Carry15a(Carry15a), .Carry15b(Carry15b), .Carry3(Carry3),
        .Carry3a(Carry3a), .Cin(Ci), .Co0_Ci0(Co0_Ci0), .Co0_Ci1(Co0_Ci1),
        .Co10_C90(Co10_C90), .Co10_C91(Co10_C91), .Co12_C110(Co12_C110),
        .Co12_C111(Co12_C111), .Co13_C120(Co13_C120), .Co13_C121(Co13_C121),
        .Co14_C130(Co14_C130), .Co14_C131(Co14_C131), .Co16_C150(Co16_C150),
        .Co16_C151(Co16_C151), .Co17_C160(Co17_C160), .Co17_C161(Co17_C161),
        .Co18_C170(Co18_C170), .Co18_C171(Co18_C171), .Co1_C00(Co1_C00),
        .Co1_C01(Co1_C01), .Co20_C190(Co20_C190), .Co20_C191(Co20_C191),
        .Co21_C200(Co21_C200), .Co21_C201(Co21_C201), .Co22_C210(Co22_C210),
        .Co22_C211(Co22_C211), .Co24_C230(Co24_C230), .Co24_C231(Co24_C231),
        .Co25_C240(Co25_C240), .Co25_C241(Co25_C241), .Co26_C250(Co26_C250),
        .Co26_C251(Co26_C251), .Co28_C270(Co28_C270), .Co28_C271(Co28_C271),
        .Co29_C280(Co29_C280), .Co29_C281(Co29_C281), .Co2_C10(Co2_C10),
        .Co2_C11(Co2_C11), .Co30_C290(Co30_C290), .Co30_C291(Co30_C291),
        .Co3_C20(Co3_C20), .Co3_C21(Co3_C21), .Co4_C30(Co4_C30),
        .Co4_C31(Co4_C31), .Co5_C40(Co5_C40), .Co5_C41(Co5_C41),
        .Co6_C50(Co6_C50), .Co6_C51(Co6_C51), .Co8_C70(Co8_C70),
        .Co8_C71(Co8_C71), .Co9_C80(Co9_C80), .Co9_C81(Co9_C81),
        .S({ S[31:0] }), .Sumi({ Sum[31:0] }) );

endmodule // add32p2

`endif

`ifdef add16p2
`else
`define add16p2
module add16p2( A , B, Ci, Co, Sum );
 input [15:0] A;
 input [15:0] B;
input Ci;
output Co;
 output [15:0] Sum;
wire [15:0] S;
wire Co6_C51;
wire Co6_C50;
wire Co5_C41;
wire Co5_C40;
wire Co4_C31;
wire Co4_C30;
wire Co3_C21;
wire Co3_C20;
wire Co2_C11;
wire Co2_C10;
wire Co1_C01;
wire Co1_C00;
wire Co0_Ci1;
wire Co0_Ci0;
wire C7_C30;
wire C7_C31;
wire Carry3;
wire C11_C70;
wire C11_C71;
wire Co8_C70;
wire Co8_C71;
wire Co9_C80;
wire Co9_C81;
wire Co10_C90;
wire Co10_C91;
wire CO12_C110;
wire Co12_C111;
wire CO13_C120;
wire Co13_C121;
wire Co14_C130;
wire Co14_C131;

sum16 I_4 ( .a({ A[0] }), .b({ B[0] }), .C11_C70(C11_C70), .C11_C71(C11_C71),
         .C7_C30(C7_C30), .C7_C31(C7_C31), .Carry3(Carry3), .Cin(Ci),
         .Co0_Ci0(Co0_Ci0), .Co0_Ci1(Co0_Ci1), .Co10_C90(Co10_C90),
         .Co10_C91(Co10_C91), .Co12_C110(CO12_C110), .Co12_C111(Co12_C111),
         .Co13_C120(CO13_C120), .Co13_C121(Co13_C121), .Co14_C130(Co14_C130),
         .Co14_C131(Co14_C131), .Co1_C00(Co1_C00), .Co1_C01(Co1_C01),
         .Co2_C10(Co2_C10), .Co2_C11(Co2_C11), .Co3_C20(Co3_C20),
         .Co3_C21(Co3_C21), .Co4_C30(Co4_C30), .Co4_C31(Co4_C31),
         .Co5_C40(Co5_C40), .Co5_C41(Co5_C41), .Co6_C50(Co6_C50),
         .Co6_C51(Co6_C51), .Co8_C70(Co8_C70), .Co8_C71(Co8_C71),
         .Co9_C80(Co9_C80), .Co9_C81(Co9_C81), .S({ S[15:0] }),
         .Sumi({ Sum[15:0] }) );
carry16 I_5 ( .a({ A[15:0] }), .b({ B[15:0] }), .C11_C70(C11_C70),
           .C11_C71(C11_C71), .C7_C30(C7_C30), .C7_C31(C7_C31),
           .Carry3(Carry3), .Co(Co), .Co0_Ci0(Co0_Ci0), .Co0_Ci1(Co0_Ci1),
           .Co10_C90(Co10_C90), .Co10_C91(Co10_C91), .Co12_C110(CO12_C110),
           .Co12_C111(Co12_C111), .Co13_C120(CO13_C120),
           .Co13_C121(Co13_C121), .Co14_C130(Co14_C130),
           .Co14_C131(Co14_C131), .Co1_C00(Co1_C00), .Co1_C01(Co1_C01),
           .Co2_C10(Co2_C10), .Co2_C11(Co2_C11), .Co3_C20(Co3_C20),
           .Co3_C21(Co3_C21), .Co4_C30(Co4_C30), .Co4_C31(Co4_C31),
           .Co5_C40(Co5_C40), .Co5_C41(Co5_C41), .Co6_C50(Co6_C50),
           .Co6_C51(Co6_C51), .Co8_C70(Co8_C70), .Co8_C71(Co8_C71),
           .Co9_C80(Co9_C80), .Co9_C81(Co9_C81), .S({ S[15:0] }) );

endmodule // add16p2

`endif

`ifdef ucebita1
`else
`define ucebita1
module ucebita1( CLK , ENH1, ENH2, ENH3, ENH4, ENL1, ENL2, ENL3, PRE, QFB, Q );
input CLK /* synthesis syn_isclock=1 */;
input PRE /* synthesis syn_isclock=1 */;
input ENH1, ENH2, ENH3, ENH4, ENL1, ENL2, ENL3;
output Q;
input QFB;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

lcell2 I_1 ( .A1(ENH2), .A2(ENL3), .A3(ENH3), .A4(ENL2), .A5(ENH4), .A6(ENL1),
          .B1(GND), .B2(GND), .C1(QFB), .C2(GND), .D1(VCC), .D2(QFB), .E1(GND),
          .E2(GND), .F1(VCC), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND),
          .MP(GND), .MS(VCC), .NP(GND), .NS(GND), .OP(ENH1), .OS(GND), .QC(CLK),
          .QR(GND), .QS(PRE), .QZ(Q) );

endmodule // ucebita1

`endif

`ifdef ucebita0
`else
`define ucebita0
module ucebita0( CLK , CLR, ENH1, ENH2, ENH3, ENH4, ENL1, ENL2, ENL3, QFB, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input ENH1, ENH2, ENH3, ENH4, ENL1, ENL2, ENL3;
output Q;
input QFB;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

lcell2 I_1 ( .A1(ENH2), .A2(ENL3), .A3(ENH3), .A4(ENL2), .A5(ENH4), .A6(ENL1),
          .B1(GND), .B2(GND), .C1(QFB), .C2(GND), .D1(VCC), .D2(QFB), .E1(GND),
          .E2(GND), .F1(VCC), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND),
          .MP(GND), .MS(VCC), .NP(GND), .NS(GND), .OP(ENH1), .OS(GND), .QC(CLK),
          .QR(CLR), .QS(GND), .QZ(Q) );

endmodule // ucebita0

`endif

`ifdef ucebit2b
`else
`define ucebit2b
module ucebit2b( CLK , CLR, ENH1, ENH2, ENH3, ENH4, ENL1, ENL2, ENL3, QFB, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input ENH1, ENH2, ENH3, ENH4, ENL1, ENL2, ENL3;
output Q;
input QFB;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

lcell2 I_1 ( .A1(ENH2), .A2(ENL3), .A3(ENH3), .A4(ENL2), .A5(ENH4), .A6(ENL1),
          .B1(GND), .B2(GND), .C1(VCC), .C2(QFB), .D1(QFB), .D2(GND), .E1(GND),
          .E2(GND), .F1(VCC), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND),
          .MP(GND), .MS(VCC), .NP(GND), .NS(GND), .OP(ENH1), .OS(GND), .QC(CLK),
          .QR(CLR), .QS(GND), .QZ(Q) );

endmodule // ucebit2b

`endif

`ifdef ttl98
`else
`define ttl98
module ttl98( A1 , A2, A3, A4, B1, B2, B3, B4, CLOCK, SEL, QA, QB, QC, QD );
input CLOCK /* synthesis syn_isclock=1 */;
input A1, A2, A3, A4, B1, B2, B3, B4;
output QA, QB, QC, QD;
input SEL;
wire N_1;
wire N_2;
wire N_3;
wire N_4;

dff QL1 ( .CLK(CLOCK), .D(N_1), .Q(QC) );
dff QL2 ( .CLK(CLOCK), .D(N_2), .Q(QD) );
dff QL3 ( .CLK(CLOCK), .D(N_3), .Q(QB) );
dff QL4 ( .CLK(CLOCK), .D(N_4), .Q(QA) );
mux2x0 QL5 ( .A(A3), .B(B3), .Q(N_1), .S(SEL) );
mux2x0 QL6 ( .A(A4), .B(B4), .Q(N_2), .S(SEL) );
mux2x0 QL7 ( .A(A2), .B(B2), .Q(N_3), .S(SEL) );
mux2x0 QL8 ( .A(A1), .B(B1), .Q(N_4), .S(SEL) );

endmodule // ttl98

`endif

`ifdef ttl91
`else
`define ttl91
module ttl91( A , B, CLK, QH, QHNN );
input CLK /* synthesis syn_isclock=1 */;
input A, B;
output QH, QHNN;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;

and2i0 QL1 ( .A(A), .B(B), .Q(N_1) );
inv QL2 ( .A(N_9), .Q(N_2) );
dff QL3 ( .CLK(CLK), .D(N_2), .Q(QHNN) );
dff QL4 ( .CLK(CLK), .D(N_9), .Q(QH) );
dff QL5 ( .CLK(CLK), .D(N_7), .Q(N_8) );
dff QL6 ( .CLK(CLK), .D(N_8), .Q(N_9) );
dff QL7 ( .CLK(CLK), .D(N_6), .Q(N_7) );
dff QL8 ( .CLK(CLK), .D(N_5), .Q(N_6) );
dff QL9 ( .CLK(CLK), .D(N_3), .Q(N_4) );
dff QL10 ( .CLK(CLK), .D(N_4), .Q(N_5) );
dff QL11 ( .CLK(CLK), .D(N_1), .Q(N_3) );

endmodule // ttl91

`endif

`ifdef ttl87
`else
`define ttl87
module ttl87( A1 , A2, A3, A4, BNN, C, Y1, Y2, Y3, Y4 );
input A1, A2, A3, A4, BNN, C;
output Y1, Y2, Y3, Y4;
wire N_1;
wire N_2;
wire N_3;
wire N_4;

and2i1 QL1 ( .A(A1), .B(BNN), .Q(N_4) );
and2i1 QL2 ( .A(A4), .B(BNN), .Q(N_1) );
and2i1 QL3 ( .A(A2), .B(BNN), .Q(N_3) );
and2i1 QL4 ( .A(A3), .B(BNN), .Q(N_2) );
xnor2i0 QL5 ( .A(N_2), .B(C), .Q(Y3) );
xnor2i0 QL6 ( .A(N_3), .B(C), .Q(Y2) );
xnor2i0 QL7 ( .A(N_4), .B(C), .Q(Y1) );
xnor2i0 QL8 ( .A(N_1), .B(C), .Q(Y4) );

endmodule // ttl87

`endif

`ifdef ttl86
`else
`define ttl86
module ttl86( A1 , A2, A3, A4, B1, B2, B3, B4, Y1, Y2, Y3, Y4 );
input A1, A2, A3, A4, B1, B2, B3, B4;
output Y1, Y2, Y3, Y4;

xor2i0 QL1 ( .A(A3), .B(B3), .Q(Y3) );
xor2i0 QL2 ( .A(A4), .B(B4), .Q(Y4) );
xor2i0 QL3 ( .A(A2), .B(B2), .Q(Y2) );
xor2i0 QL4 ( .A(A1), .B(B1), .Q(Y1) );

endmodule // ttl86

`endif

`ifdef ttl85
`else
`define ttl85
module ttl85( A0 , A1, A2, A3, AEQB, AGTB, ALTB, B0, B1, B2, B3, AEQBO, AGTBO,
              ALTBO );
input A0, A1, A2, A3, AEQB;
output AEQBO;
input AGTB;
output AGTBO;
input ALTB;
output ALTBO;
input B0, B1, B2, B3;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;
wire N_15;
wire N_16;
wire N_17;
wire N_18;
wire N_19;
wire N_20;
wire N_21;
wire N_22;
wire N_23;

and2i1 QL26 ( .A(B3), .B(A3), .Q(N_4) );
and2i1 QL25 ( .A(A3), .B(B3), .Q(N_3) );
and2i1 QL24 ( .A(B0), .B(A0), .Q(N_6) );
and2i1 QL23 ( .A(A0), .B(B0), .Q(N_5) );
and2i1 QL22 ( .A(A2), .B(B2), .Q(N_7) );
and2i1 QL21 ( .A(B2), .B(A2), .Q(N_8) );
and2i1 QL20 ( .A(A3), .B(B3), .Q(N_17) );
and2i1 QL19 ( .A(B1), .B(A1), .Q(N_10) );
and2i1 QL18 ( .A(A1), .B(B1), .Q(N_9) );
and2i1 QL17 ( .A(B3), .B(A3), .Q(N_23) );
or2i0 QL16 ( .A(N_6), .B(N_5), .Q(N_11) );
or2i0 QL15 ( .A(N_10), .B(N_9), .Q(N_12) );
nor2i0 QL14 ( .A(N_4), .B(N_3), .Q(N_1) );
nor2i0 QL13 ( .A(N_8), .B(N_7), .Q(N_2) );
and3i1 QL12 ( .A(N_1), .B(B2), .C(A2), .Q(N_16) );
and3i1 QL11 ( .A(N_1), .B(A2), .C(B2), .Q(N_15) );
and4i1 QL10 ( .A(N_1), .B(N_2), .C(B1), .D(A1), .Q(N_14) );
and4i1 QL9 ( .A(N_1), .B(N_2), .C(A1), .D(B1), .Q(N_18) );
and5i2 QL8 ( .A(N_1), .B(N_2), .C(B0), .D(N_12), .E(A0), .Q(N_19) );
and5i2 QL7 ( .A(N_1), .B(N_2), .C(A0), .D(N_12), .E(B0), .Q(N_20) );
and5i2 QL6 ( .A(N_1), .B(N_2), .C(AGTB), .D(N_12), .E(N_11), .Q(N_21) );
and5i2 QL5 ( .A(N_1), .B(N_2), .C(ALTB), .D(N_12), .E(N_11), .Q(N_13) );
and5i2 QL4 ( .A(N_1), .B(N_2), .C(AEQB), .D(N_12), .E(N_11), .Q(AEQBO) );
or5i0 QL3 ( .A(N_22), .B(N_16), .C(N_14), .D(N_19), .E(N_13), .Q(ALTBO) );
or5i0 QL2 ( .A(N_17), .B(N_15), .C(N_18), .D(N_20), .E(N_21), .Q(AGTBO) );
buff QL1 ( .A(N_23), .Q(N_22) );

endmodule // ttl85

`endif

`ifdef ttl842q
`else
`define ttl842q
module ttl842q( D1 , D10, D2, D3, D4, D5, D6, D7, D8, D9, G, Q1, Q10, Q2, Q3, Q4,
                Q5, Q6, Q7, Q8, Q9 );
input D1, D10, D2, D3, D4, D5, D6, D7, D8, D9, G;
output Q1, Q10, Q2, Q3, Q4, Q5, Q6, Q7, Q8, Q9;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;

inv QL1 ( .A(D10), .Q(N_8) );
inv QL2 ( .A(D9), .Q(N_1) );
inv QL3 ( .A(D8), .Q(N_9) );
inv QL4 ( .A(D7), .Q(N_2) );
inv QL5 ( .A(D6), .Q(N_10) );
inv QL6 ( .A(D5), .Q(N_3) );
inv QL7 ( .A(D4), .Q(N_5) );
inv QL8 ( .A(D3), .Q(N_4) );
inv QL9 ( .A(D2), .Q(N_7) );
inv QL10 ( .A(D1), .Q(N_6) );
dlad QL11 ( .D1(N_1), .D2(N_8), .G(G), .Q1(Q9), .Q2(Q10) );
dlad QL12 ( .D1(N_2), .D2(N_9), .G(G), .Q1(Q7), .Q2(Q8) );
dlad QL13 ( .D1(N_3), .D2(N_10), .G(G), .Q1(Q5), .Q2(Q6) );
dlad QL14 ( .D1(N_4), .D2(N_5), .G(G), .Q1(Q3), .Q2(Q4) );
dlad QL15 ( .D1(N_6), .D2(N_7), .G(G), .Q1(Q1), .Q2(Q2) );

endmodule // ttl842q

`endif

`ifdef ttl841q
`else
`define ttl841q
module ttl841q( D1 , D10, D2, D3, D4, D5, D6, D7, D8, D9, G, Q1, Q10, Q2, Q3, Q4,
                Q5, Q6, Q7, Q8, Q9 );
input D1, D10, D2, D3, D4, D5, D6, D7, D8, D9, G;
output Q1, Q10, Q2, Q3, Q4, Q5, Q6, Q7, Q8, Q9;

dlad QL1 ( .D1(D9), .D2(D10), .G(G), .Q1(Q9), .Q2(Q10) );
dlad QL2 ( .D1(D7), .D2(D8), .G(G), .Q1(Q7), .Q2(Q8) );
dlad QL3 ( .D1(D5), .D2(D6), .G(G), .Q1(Q5), .Q2(Q6) );
dlad QL4 ( .D1(D3), .D2(D4), .G(G), .Q1(Q3), .Q2(Q4) );
dlad QL5 ( .D1(D1), .D2(D2), .G(G), .Q1(Q1), .Q2(Q2) );

endmodule // ttl841q

`endif

`ifdef ttl823q
`else
`define ttl823q
module ttl823q( CLK , CLKENBLNN, CLR, D1, D2, D3, D4, D5, D6, D7, D8, D9, Q1, Q2,
                Q3, Q4, Q5, Q6, Q7, Q8, Q9 );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input CLKENBLNN, D1, D2, D3, D4, D5, D6, D7, D8, D9;
output Q1, Q2, Q3, Q4, Q5, Q6, Q7, Q8, Q9;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;

dffc QL1 ( .CLK(CLK), .CLR(CLR), .D(N_1), .Q(Q9) );
dffc QL2 ( .CLK(CLK), .CLR(CLR), .D(N_2), .Q(Q8) );
dffc QL3 ( .CLK(CLK), .CLR(CLR), .D(N_9), .Q(Q7) );
dffc QL4 ( .CLK(CLK), .CLR(CLR), .D(N_8), .Q(Q6) );
dffc QL5 ( .CLK(CLK), .CLR(CLR), .D(N_7), .Q(Q5) );
dffc QL6 ( .CLK(CLK), .CLR(CLR), .D(N_6), .Q(Q4) );
dffc QL7 ( .CLK(CLK), .CLR(CLR), .D(N_5), .Q(Q3) );
dffc QL8 ( .CLK(CLK), .CLR(CLR), .D(N_4), .Q(Q2) );
dffc QL9 ( .CLK(CLK), .CLR(CLR), .D(N_3), .Q(Q1) );
mux2x0 QL10 ( .A(D9), .B(Q9), .Q(N_1), .S(CLKENBLNN) );
mux2x0 QL11 ( .A(D8), .B(Q8), .Q(N_2), .S(CLKENBLNN) );
mux2x0 QL12 ( .A(D7), .B(Q7), .Q(N_9), .S(CLKENBLNN) );
mux2x0 QL13 ( .A(D6), .B(Q6), .Q(N_8), .S(CLKENBLNN) );
mux2x0 QL14 ( .A(D5), .B(Q5), .Q(N_7), .S(CLKENBLNN) );
mux2x0 QL15 ( .A(D4), .B(Q4), .Q(N_6), .S(CLKENBLNN) );
mux2x0 QL16 ( .A(D3), .B(Q3), .Q(N_5), .S(CLKENBLNN) );
mux2x0 QL17 ( .A(D2), .B(Q2), .Q(N_4), .S(CLKENBLNN) );
mux2x0 QL18 ( .A(D1), .B(Q1), .Q(N_3), .S(CLKENBLNN) );

endmodule // ttl823q

`endif

`ifdef ttl822
`else
`define ttl822
module ttl822( CLK , D1, D10, D2, D3, D4, D5, D6, D7, D8, D9, Q1, Q10, Q2, Q3, Q4,
               Q5, Q6, Q7, Q8, Q9 );
input CLK /* synthesis syn_isclock=1 */;
input D1, D10, D2, D3, D4, D5, D6, D7, D8, D9;
output Q1, Q10, Q2, Q3, Q4, Q5, Q6, Q7, Q8, Q9;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;

inv QL1 ( .A(D10), .Q(N_1) );
inv QL2 ( .A(D9), .Q(N_2) );
inv QL3 ( .A(D8), .Q(N_3) );
inv QL4 ( .A(D7), .Q(N_4) );
inv QL5 ( .A(D6), .Q(N_5) );
inv QL6 ( .A(D5), .Q(N_6) );
inv QL7 ( .A(D4), .Q(N_7) );
inv QL8 ( .A(D3), .Q(N_8) );
inv QL9 ( .A(D2), .Q(N_9) );
inv QL10 ( .A(D1), .Q(N_10) );
dff QL11 ( .CLK(CLK), .D(N_1), .Q(Q10) );
dff QL12 ( .CLK(CLK), .D(N_2), .Q(Q9) );
dff QL13 ( .CLK(CLK), .D(N_3), .Q(Q8) );
dff QL14 ( .CLK(CLK), .D(N_4), .Q(Q7) );
dff QL15 ( .CLK(CLK), .D(N_5), .Q(Q6) );
dff QL16 ( .CLK(CLK), .D(N_6), .Q(Q5) );
dff QL17 ( .CLK(CLK), .D(N_7), .Q(Q4) );
dff QL18 ( .CLK(CLK), .D(N_8), .Q(Q3) );
dff QL19 ( .CLK(CLK), .D(N_9), .Q(Q2) );
dff QL20 ( .CLK(CLK), .D(N_10), .Q(Q1) );

endmodule // ttl822

`endif

`ifdef ttl821
`else
`define ttl821
module ttl821( CLK , D1, D10, D2, D3, D4, D5, D6, D7, D8, D9, Q1, Q10, Q2, Q3, Q4,
               Q5, Q6, Q7, Q8, Q9 );
input CLK /* synthesis syn_isclock=1 */;
input D1, D10, D2, D3, D4, D5, D6, D7, D8, D9;
output Q1, Q10, Q2, Q3, Q4, Q5, Q6, Q7, Q8, Q9;

dff QL1 ( .CLK(CLK), .D(D10), .Q(Q10) );
dff QL2 ( .CLK(CLK), .D(D9), .Q(Q9) );
dff QL3 ( .CLK(CLK), .D(D8), .Q(Q8) );
dff QL4 ( .CLK(CLK), .D(D7), .Q(Q7) );
dff QL5 ( .CLK(CLK), .D(D6), .Q(Q6) );
dff QL6 ( .CLK(CLK), .D(D5), .Q(Q5) );
dff QL7 ( .CLK(CLK), .D(D4), .Q(Q4) );
dff QL8 ( .CLK(CLK), .D(D3), .Q(Q3) );
dff QL9 ( .CLK(CLK), .D(D2), .Q(Q2) );
dff QL10 ( .CLK(CLK), .D(D1), .Q(Q1) );

endmodule // ttl821

`endif

`ifdef ttl78q
`else
`define ttl78q
module ttl78q( CLK , CLR, J1, J2, K1, K2, PRE1, PRE2, Q1, Q2 );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input PRE1 /* synthesis syn_isclock=1 */;
input PRE2 /* synthesis syn_isclock=1 */;
input J1, J2, K1, K2;
output Q1, Q2;

jkffpc QL1 ( .CLK(CLK), .CLR(CLR), .J(J2), .K(K2), .PRE(PRE2), .Q(Q2) );
jkffpc QL2 ( .CLK(CLK), .CLR(CLR), .J(J1), .K(K1), .PRE(PRE1), .Q(Q1) );

endmodule // ttl78q

`endif

`ifdef ttl77
`else
`define ttl77
module ttl77( C1C2 , C3C4, D1, D2, D3, D4, Q1, Q2, Q3, Q4 );
input C1C2, C3C4, D1, D2, D3, D4;
output Q1, Q2, Q3, Q4;

dlad QL1 ( .D1(D3), .D2(D4), .G(C3C4), .Q1(Q3), .Q2(Q4) );
dlad QL2 ( .D1(D1), .D2(D2), .G(C1C2), .Q1(Q1), .Q2(Q2) );

endmodule // ttl77

`endif

`ifdef ttl74q
`else
`define ttl74q
module ttl74q( CLK1 , CLK2, CLR1, CLR2, D1, D2, PRE1, PRE2, Q1, Q2 );
input CLK1 /* synthesis syn_isclock=1 */;
input CLK2 /* synthesis syn_isclock=1 */;
input CLR1 /* synthesis syn_isclock=1 */;
input CLR2 /* synthesis syn_isclock=1 */;
input PRE1 /* synthesis syn_isclock=1 */;
input PRE2 /* synthesis syn_isclock=1 */;
input D1, D2;
output Q1, Q2;

dffpc QL1 ( .CLK(CLK2), .CLR(CLR2), .D(D2), .PRE(PRE2), .Q(Q2) );
dffpc QL2 ( .CLK(CLK1), .CLR(CLR1), .D(D1), .PRE(PRE1), .Q(Q1) );

endmodule // ttl74q

`endif

`ifdef ttl688
`else
`define ttl688
module ttl688( GNN , P0, P1, P2, P3, P4, P5, P6, P7, Q0, Q1, Q2, Q3, Q4, Q5, Q6,
               Q7, PQ );
input GNN, P0, P1, P2, P3, P4, P5, P6, P7;
output PQ;
input Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7;
supply0 GND;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;

nand13i6 QL1 ( .A(N_1), .B(N_2), .C(N_3), .D(N_4), .E(N_5), .F(N_6), .G(N_7),
            .H(N_8), .I(GNN), .J(GND), .K(GND), .L(GND), .M(GND), .Q(PQ) );
xnor2i0 QL2 ( .A(Q1), .B(P1), .Q(N_7) );
xnor2i0 QL3 ( .A(Q2), .B(P2), .Q(N_6) );
xnor2i0 QL4 ( .A(Q7), .B(P7), .Q(N_1) );
xnor2i0 QL5 ( .A(Q6), .B(P6), .Q(N_2) );
xnor2i0 QL6 ( .A(Q5), .B(P5), .Q(N_3) );
xnor2i0 QL7 ( .A(Q4), .B(P4), .Q(N_4) );
xnor2i0 QL8 ( .A(Q3), .B(P3), .Q(N_5) );
xor2i0 QL9 ( .A(Q0), .B(P0), .Q(N_8) );

endmodule // ttl688

`endif

`ifdef ttl686
`else
`define ttl686
module ttl686( G1NN , G2NN, P0, P1, P2, P3, P4, P5, P6, P7, Q0, Q1, Q2, Q3, Q4, Q5,
               Q6, Q7, PGTRQ, PQ );
input G1NN, G2NN, P0, P1, P2, P3, P4, P5, P6, P7;
output PGTRQ, PQ;
input Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
supply1 VCC;
supply0 GND;
wire N_11;
wire N_12;
wire N_13;
wire N_14;
wire N_15;
wire N_16;
wire N_17;

and3i2 QL1 ( .A(P6), .B(N_17), .C(Q6), .Q(N_3) );
and4i3 QL2 ( .A(P5), .B(N_17), .C(N_16), .D(Q5), .Q(N_9) );
and5i4 QL3 ( .A(P4), .B(N_17), .C(N_16), .D(N_15), .E(Q4), .Q(N_8) );
and6i5 QL4 ( .A(P3), .B(N_17), .C(N_16), .D(N_15), .E(N_10), .F(Q3), .Q(N_7) );
nand2i1 QL5 ( .A(P7), .B(Q7), .Q(N_2) );
or2i0 QL6 ( .A(G2NN), .B(N_1), .Q(PGTRQ) );
xnor2i0 QL7 ( .A(Q0), .B(P0), .Q(N_11) );
xnor2i0 QL8 ( .A(Q1), .B(P1), .Q(N_12) );
xnor2i0 QL9 ( .A(Q3), .B(P3), .Q(N_14) );
xnor2i0 QL10 ( .A(Q2), .B(P2), .Q(N_13) );
and14i7 QL11 ( .A(VCC), .B(VCC), .C(VCC), .D(VCC), .E(VCC), .F(VCC), .G(N_2),
            .H(N_4), .I(N_5), .J(N_6), .K(N_7), .L(N_8), .M(N_9), .N(N_3),
            .Q(N_1) );
and14i7 QL12 ( .A(P2), .B(VCC), .C(VCC), .D(VCC), .E(VCC), .F(VCC), .G(N_14),
            .H(N_10), .I(Q2), .J(N_15), .K(N_16), .L(N_17), .M(GND), .N(GND),
            .Q(N_6) );
and14i7 QL13 ( .A(P1), .B(VCC), .C(VCC), .D(N_13), .E(N_14), .F(VCC), .G(VCC),
            .H(N_10), .I(N_15), .J(Q1), .K(N_16), .L(N_17), .M(GND), .N(GND),
            .Q(N_5) );
and14i7 QL14 ( .A(P0), .B(VCC), .C(VCC), .D(N_12), .E(N_13), .F(N_14), .G(VCC),
            .H(N_10), .I(N_15), .J(N_16), .K(Q0), .L(N_17), .M(GND), .N(GND),
            .Q(N_4) );
xor2i0 QL15 ( .A(Q7), .B(P7), .Q(N_17) );
xor2i0 QL16 ( .A(Q6), .B(P6), .Q(N_16) );
xor2i0 QL17 ( .A(Q5), .B(P5), .Q(N_15) );
xor2i0 QL18 ( .A(Q4), .B(P4), .Q(N_10) );
or13i6 QL19 ( .A(N_17), .B(N_16), .C(N_15), .D(N_10), .E(GND), .F(G1NN), .G(GND),
           .H(N_14), .I(N_13), .J(N_12), .K(N_11), .L(VCC), .M(VCC), .Q(PQ) );

endmodule // ttl686

`endif

`ifdef ttl684
`else
`define ttl684
module ttl684( P0 , P1, P2, P3, P4, P5, P6, P7, Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7,
               PGTRQ, PQ );
input P0, P1, P2, P3, P4, P5, P6, P7;
output PGTRQ, PQ;
input Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
supply1 VCC;
supply0 GND;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;
wire N_15;
wire N_16;

and3i2 QL1 ( .A(P6), .B(N_16), .C(Q6), .Q(N_2) );
and4i3 QL2 ( .A(P5), .B(N_16), .C(N_15), .D(Q5), .Q(N_8) );
and5i4 QL3 ( .A(P4), .B(N_16), .C(N_15), .D(N_14), .E(Q4), .Q(N_7) );
and6i5 QL4 ( .A(P3), .B(N_16), .C(N_15), .D(N_14), .E(N_9), .F(Q3), .Q(N_6) );
nand2i1 QL5 ( .A(P7), .B(Q7), .Q(N_1) );
xnor2i0 QL6 ( .A(Q0), .B(P0), .Q(N_10) );
xnor2i0 QL7 ( .A(Q1), .B(P1), .Q(N_11) );
xnor2i0 QL8 ( .A(Q3), .B(P3), .Q(N_13) );
xnor2i0 QL9 ( .A(Q2), .B(P2), .Q(N_12) );
and14i7 QL10 ( .A(VCC), .B(VCC), .C(VCC), .D(VCC), .E(VCC), .F(VCC), .G(N_1),
            .H(N_3), .I(N_4), .J(N_5), .K(N_6), .L(N_7), .M(N_8), .N(N_2),
            .Q(PGTRQ) );
and14i7 QL11 ( .A(P2), .B(VCC), .C(VCC), .D(VCC), .E(VCC), .F(VCC), .G(N_13),
            .H(N_9), .I(Q2), .J(N_14), .K(N_15), .L(N_16), .M(GND), .N(GND),
            .Q(N_5) );
and14i7 QL12 ( .A(P1), .B(VCC), .C(VCC), .D(N_12), .E(N_13), .F(VCC), .G(VCC),
            .H(N_9), .I(N_14), .J(Q1), .K(N_15), .L(N_16), .M(GND), .N(GND),
            .Q(N_4) );
and14i7 QL13 ( .A(P0), .B(VCC), .C(VCC), .D(N_11), .E(N_12), .F(N_13), .G(VCC),
            .H(N_9), .I(N_14), .J(N_15), .K(Q0), .L(N_16), .M(GND), .N(GND),
            .Q(N_3) );
xor2i0 QL14 ( .A(Q7), .B(P7), .Q(N_16) );
xor2i0 QL15 ( .A(Q6), .B(P6), .Q(N_15) );
xor2i0 QL16 ( .A(Q5), .B(P5), .Q(N_14) );
xor2i0 QL17 ( .A(Q4), .B(P4), .Q(N_9) );
or13i6 QL18 ( .A(N_16), .B(N_15), .C(N_14), .D(N_9), .E(GND), .F(GND), .G(GND),
           .H(N_13), .I(N_12), .J(N_11), .K(N_10), .L(VCC), .M(VCC), .Q(PQ) );

endmodule // ttl684

`endif

`ifdef ttl604q
`else
`define ttl604q
module ttl604q( A1 , A2, A3, A4, A5, A6, A7, A8, B1, B2, B3, B4, B5, B6, B7, B8,
                CLK, SEL, Y1, Y2, Y3, Y4, Y5, Y6, Y7, Y8 );
input A1, A2, A3, A4, A5, A6, A7, A8, B1, B2, B3, B4, B5, B6, B7, B8, CLK,
SEL;
output Y1, Y2, Y3, Y4, Y5, Y6, Y7, Y8;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;
wire N_15;
wire N_16;

mux2x0 QL1 ( .A(N_16), .B(N_8), .Q(Y8), .S(SEL) );
mux2x0 QL2 ( .A(N_15), .B(N_7), .Q(Y7), .S(SEL) );
mux2x0 QL3 ( .A(N_14), .B(N_6), .Q(Y6), .S(SEL) );
mux2x0 QL4 ( .A(N_13), .B(N_5), .Q(Y5), .S(SEL) );
mux2x0 QL5 ( .A(N_9), .B(N_1), .Q(Y1), .S(SEL) );
mux2x0 QL6 ( .A(N_12), .B(N_4), .Q(Y4), .S(SEL) );
mux2x0 QL7 ( .A(N_11), .B(N_3), .Q(Y3), .S(SEL) );
mux2x0 QL8 ( .A(N_10), .B(N_2), .Q(Y2), .S(SEL) );
dff QL9 ( .CLK(CLK), .D(B8), .Q(N_16) );
dff QL10 ( .CLK(CLK), .D(A8), .Q(N_8) );
dff QL11 ( .CLK(CLK), .D(B7), .Q(N_15) );
dff QL12 ( .CLK(CLK), .D(A7), .Q(N_7) );
dff QL13 ( .CLK(CLK), .D(B6), .Q(N_14) );
dff QL14 ( .CLK(CLK), .D(A6), .Q(N_6) );
dff QL15 ( .CLK(CLK), .D(B5), .Q(N_13) );
dff QL16 ( .CLK(CLK), .D(A5), .Q(N_5) );
dff QL17 ( .CLK(CLK), .D(B1), .Q(N_9) );
dff QL18 ( .CLK(CLK), .D(A1), .Q(N_1) );
dff QL19 ( .CLK(CLK), .D(B4), .Q(N_12) );
dff QL20 ( .CLK(CLK), .D(A4), .Q(N_4) );
dff QL21 ( .CLK(CLK), .D(B3), .Q(N_11) );
dff QL22 ( .CLK(CLK), .D(A3), .Q(N_3) );
dff QL23 ( .CLK(CLK), .D(B2), .Q(N_10) );
dff QL24 ( .CLK(CLK), .D(A2), .Q(N_2) );

endmodule // ttl604q

`endif

`ifdef ttl595q
`else
`define ttl595q
module ttl595q( RCLK , SER, SRCLK, SRCLR, QA, QB, QC, QD, QE, QF, QG, QH, QHNN );
output QA, QB, QC, QD, QE, QF, QG, QH, QHNN;
input RCLK /* synthesis syn_isclock=1 */;
input SRCLK /* synthesis syn_isclock=1 */;
input SRCLR /* synthesis syn_isclock=1 */;
input SER;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;

inv QL1 ( .A(QHNN), .Q(N_1) );
inv QL2 ( .A(N_3), .Q(N_2) );
dffp QL3 ( .CLK(SRCLK), .D(N_2), .PRE(SRCLR), .Q(QHNN) );
dff QL4 ( .CLK(RCLK), .D(N_1), .Q(QH) );
dff QL5 ( .CLK(RCLK), .D(N_3), .Q(QG) );
dff QL6 ( .CLK(RCLK), .D(N_9), .Q(QF) );
dff QL7 ( .CLK(RCLK), .D(N_8), .Q(QE) );
dff QL8 ( .CLK(RCLK), .D(N_7), .Q(QD) );
dff QL9 ( .CLK(RCLK), .D(N_6), .Q(QC) );
dff QL10 ( .CLK(RCLK), .D(N_5), .Q(QB) );
dff QL11 ( .CLK(RCLK), .D(N_4), .Q(QA) );
dffc QL12 ( .CLK(SRCLK), .CLR(SRCLR), .D(N_9), .Q(N_3) );
dffc QL13 ( .CLK(SRCLK), .CLR(SRCLR), .D(N_8), .Q(N_9) );
dffc QL14 ( .CLK(SRCLK), .CLR(SRCLR), .D(N_7), .Q(N_8) );
dffc QL15 ( .CLK(SRCLK), .CLR(SRCLR), .D(N_6), .Q(N_7) );
dffc QL16 ( .CLK(SRCLK), .CLR(SRCLR), .D(N_5), .Q(N_6) );
dffc QL17 ( .CLK(SRCLK), .CLR(SRCLR), .D(N_4), .Q(N_5) );
dffc QL18 ( .CLK(SRCLK), .CLR(SRCLR), .D(SER), .Q(N_4) );

endmodule // ttl595q

`endif

`ifdef ttl594q
`else
`define ttl594q
module ttl594q( RCLK , RCLR, SER, SRCLK, SRCLR, QA, QB, QC, QD, QE, QF, QG, QH,
                QHNN );
output QA, QB, QC, QD, QE, QF, QG, QH, QHNN;
input RCLK /* synthesis syn_isclock=1 */;
input RCLR /* synthesis syn_isclock=1 */;
input SRCLK /* synthesis syn_isclock=1 */;
input SRCLR /* synthesis syn_isclock=1 */;
input SER;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;

inv QL1 ( .A(QHNN), .Q(N_1) );
inv QL2 ( .A(N_3), .Q(N_2) );
dffp QL3 ( .CLK(SRCLK), .D(N_2), .PRE(SRCLR), .Q(QHNN) );
dffc QL4 ( .CLK(RCLK), .CLR(RCLR), .D(N_1), .Q(QH) );
dffc QL5 ( .CLK(RCLK), .CLR(RCLR), .D(N_3), .Q(QG) );
dffc QL6 ( .CLK(RCLK), .CLR(RCLR), .D(N_4), .Q(QA) );
dffc QL7 ( .CLK(RCLK), .CLR(RCLR), .D(N_6), .Q(QC) );
dffc QL8 ( .CLK(RCLK), .CLR(RCLR), .D(N_8), .Q(QE) );
dffc QL9 ( .CLK(RCLK), .CLR(RCLR), .D(N_7), .Q(QD) );
dffc QL10 ( .CLK(RCLK), .CLR(RCLR), .D(N_9), .Q(QF) );
dffc QL11 ( .CLK(RCLK), .CLR(RCLR), .D(N_5), .Q(QB) );
dffc QL12 ( .CLK(SRCLK), .CLR(SRCLR), .D(N_9), .Q(N_3) );
dffc QL13 ( .CLK(SRCLK), .CLR(SRCLR), .D(N_8), .Q(N_9) );
dffc QL14 ( .CLK(SRCLK), .CLR(SRCLR), .D(N_7), .Q(N_8) );
dffc QL15 ( .CLK(SRCLK), .CLR(SRCLR), .D(N_6), .Q(N_7) );
dffc QL16 ( .CLK(SRCLK), .CLR(SRCLR), .D(N_5), .Q(N_6) );
dffc QL17 ( .CLK(SRCLK), .CLR(SRCLR), .D(N_4), .Q(N_5) );
dffc QL18 ( .CLK(SRCLK), .CLR(SRCLR), .D(SER), .Q(N_4) );

endmodule // ttl594q

`endif

`ifdef ttl518
`else
`define ttl518
module ttl518( GNN , P0, P1, P2, P3, P4, P5, P6, P7, Q0, Q1, Q2, Q3, Q4, Q5, Q6,
               Q7, PQ );
input GNN, P0, P1, P2, P3, P4, P5, P6, P7;
output PQ;
input Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7;
supply0 GND;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;

xnor2i0 QL1 ( .A(Q7), .B(P7), .Q(N_1) );
xnor2i0 QL2 ( .A(Q6), .B(P6), .Q(N_2) );
xnor2i0 QL3 ( .A(Q5), .B(P5), .Q(N_3) );
xnor2i0 QL4 ( .A(Q4), .B(P4), .Q(N_4) );
xnor2i0 QL5 ( .A(Q3), .B(P3), .Q(N_5) );
xnor2i0 QL6 ( .A(Q2), .B(P2), .Q(N_6) );
xnor2i0 QL7 ( .A(Q1), .B(P1), .Q(N_7) );
and14i7 QL8 ( .A(N_1), .B(N_2), .C(N_3), .D(N_4), .E(N_5), .F(N_6), .G(N_7), .H(N_8),
           .I(GNN), .J(GND), .K(GND), .L(GND), .M(GND), .N(GND), .Q(PQ) );
xor2i0 QL9 ( .A(Q0), .B(P0), .Q(N_8) );

endmodule // ttl518

`endif

`ifdef ttl468
`else
`define ttl468
module ttl468( A1_1 , A1_2, A1_3, A1_4, A2_1, A2_2, A2_3, A2_4, G1NN, G2NN, Y1_1,
               Y1_2, Y1_3, Y1_4, Y2_1, Y2_2, Y2_3, Y2_4 );
input A1_1, A1_2, A1_3, A1_4, A2_1, A2_2, A2_3, A2_4, G1NN, G2NN;
output Y1_1, Y1_2, Y1_3, Y1_4, Y2_1, Y2_2, Y2_3, Y2_4;
wire N_1;
wire N_2;

inv QL1 ( .A(G2NN), .Q(N_2) );
inv QL2 ( .A(G1NN), .Q(N_1) );
triipad QL3 ( .A(A2_4), .EN(N_2), .P(Y2_4) );
triipad QL4 ( .A(A2_3), .EN(N_2), .P(Y2_3) );
triipad QL5 ( .A(A2_2), .EN(N_2), .P(Y2_2) );
triipad QL6 ( .A(A2_1), .EN(N_2), .P(Y2_1) );
triipad QL7 ( .A(A1_3), .EN(N_1), .P(Y1_3) );
triipad QL8 ( .A(A1_4), .EN(N_1), .P(Y1_4) );
triipad QL9 ( .A(A1_2), .EN(N_1), .P(Y1_2) );
triipad QL10 ( .A(A1_1), .EN(N_1), .P(Y1_1) );

endmodule // ttl468

`endif

`ifdef ttl467
`else
`define ttl467
module ttl467( A1_1 , A1_2, A1_3, A1_4, A2_1, A2_2, A2_3, A2_4, G1NN, G2NN, Y1_1,
               Y1_2, Y1_3, Y1_4, Y2_1, Y2_2, Y2_3, Y2_4 );
input A1_1, A1_2, A1_3, A1_4, A2_1, A2_2, A2_3, A2_4, G1NN, G2NN;
output Y1_1, Y1_2, Y1_3, Y1_4, Y2_1, Y2_2, Y2_3, Y2_4;
wire N_1;
wire N_2;

inv QL1 ( .A(G2NN), .Q(N_2) );
inv QL2 ( .A(G1NN), .Q(N_1) );
tripad QL3 ( .A(A2_4), .EN(N_2), .P(Y2_4) );
tripad QL4 ( .A(A2_3), .EN(N_2), .P(Y2_3) );
tripad QL5 ( .A(A2_2), .EN(N_2), .P(Y2_2) );
tripad QL6 ( .A(A2_1), .EN(N_2), .P(Y2_1) );
tripad QL7 ( .A(A1_4), .EN(N_1), .P(Y1_4) );
tripad QL8 ( .A(A1_3), .EN(N_1), .P(Y1_3) );
tripad QL9 ( .A(A1_2), .EN(N_1), .P(Y1_2) );
tripad QL10 ( .A(A1_1), .EN(N_1), .P(Y1_1) );

endmodule // ttl467

`endif

`ifdef ttl466
`else
`define ttl466
module ttl466( A1 , A2, A3, A4, A5, A6, A7, A8, G1NN, G2NN, Y1, Y2, Y3, Y4, Y5,
               Y6, Y7, Y8 );
input A1, A2, A3, A4, A5, A6, A7, A8, G1NN, G2NN;
output Y1, Y2, Y3, Y4, Y5, Y6, Y7, Y8;
wire N_1;

triipad QL1 ( .A(A3), .EN(N_1), .P(Y3) );
triipad QL2 ( .A(A8), .EN(N_1), .P(Y8) );
triipad QL3 ( .A(A7), .EN(N_1), .P(Y7) );
triipad QL4 ( .A(A6), .EN(N_1), .P(Y6) );
triipad QL5 ( .A(A5), .EN(N_1), .P(Y5) );
triipad QL6 ( .A(A4), .EN(N_1), .P(Y4) );
triipad QL7 ( .A(A2), .EN(N_1), .P(Y2) );
triipad QL8 ( .A(A1), .EN(N_1), .P(Y1) );
and2i2 QL9 ( .A(G1NN), .B(G2NN), .Q(N_1) );

endmodule // ttl466

`endif

`ifdef ttl465
`else
`define ttl465
module ttl465( A1 , A2, A3, A4, A5, A6, A7, A8, G1NN, G2NN, Y1, Y2, Y3, Y4, Y5,
               Y6, Y7, Y8 );
input A1, A2, A3, A4, A5, A6, A7, A8, G1NN, G2NN;
output Y1, Y2, Y3, Y4, Y5, Y6, Y7, Y8;
wire N_1;

and2i2 QL1 ( .A(G1NN), .B(G2NN), .Q(N_1) );
tripad QL2 ( .A(A8), .EN(N_1), .P(Y8) );
tripad QL3 ( .A(A7), .EN(N_1), .P(Y7) );
tripad QL4 ( .A(A6), .EN(N_1), .P(Y6) );
tripad QL5 ( .A(A5), .EN(N_1), .P(Y5) );
tripad QL6 ( .A(A2), .EN(N_1), .P(Y2) );
tripad QL7 ( .A(A4), .EN(N_1), .P(Y4) );
tripad QL8 ( .A(A3), .EN(N_1), .P(Y3) );
tripad QL9 ( .A(A1), .EN(N_1), .P(Y1) );

endmodule // ttl465

`endif

`ifdef ttl42q
`else
`define ttl42q
module ttl42q( A , B, C, D, Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7, Q8, Q9 );
input A, B, C, D;
output Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7, Q8, Q9;

and4i4 QL1 ( .A(A), .B(B), .C(C), .D(D), .Q(Q0) );
and4i1 QL2 ( .A(A), .B(B), .C(C), .D(D), .Q(Q7) );
and4i2 QL3 ( .A(A), .B(D), .C(B), .D(C), .Q(Q9) );
and4i2 QL4 ( .A(B), .B(C), .C(A), .D(D), .Q(Q6) );
and4i2 QL5 ( .A(A), .B(C), .C(B), .D(D), .Q(Q5) );
and4i2 QL6 ( .A(A), .B(B), .C(C), .D(D), .Q(Q3) );
and4i3 QL7 ( .A(D), .B(A), .C(B), .D(C), .Q(Q8) );
and4i3 QL8 ( .A(C), .B(A), .C(B), .D(D), .Q(Q4) );
and4i3 QL9 ( .A(B), .B(A), .C(C), .D(D), .Q(Q2) );
and4i3 QL10 ( .A(A), .B(B), .C(C), .D(D), .Q(Q1) );

endmodule // ttl42q

`endif

`ifdef ttl396
`else
`define ttl396
module ttl396( CLK , D1, D2, D3, D4, GNN, Q1_1, Q1_2, Q2_1, Q2_2, Q3_1, Q3_2,
               Q4_1, Q4_2 );
input CLK /* synthesis syn_isclock=1 */;
input D1, D2, D3, D4, GNN;
output Q1_1, Q1_2, Q2_1, Q2_2, Q3_1, Q3_2, Q4_1, Q4_2;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;

and2i1 QL1 ( .A(N_4), .B(GNN), .Q(Q4_2) );
and2i1 QL2 ( .A(N_5), .B(GNN), .Q(Q4_1) );
and2i1 QL3 ( .A(N_6), .B(GNN), .Q(Q3_2) );
and2i1 QL4 ( .A(N_1), .B(GNN), .Q(Q3_1) );
and2i1 QL5 ( .A(N_7), .B(GNN), .Q(Q2_2) );
and2i1 QL6 ( .A(N_2), .B(GNN), .Q(Q1_2) );
and2i1 QL7 ( .A(N_8), .B(GNN), .Q(Q2_1) );
and2i1 QL8 ( .A(N_3), .B(GNN), .Q(Q1_1) );
dff QL9 ( .CLK(CLK), .D(N_3), .Q(N_8) );
dff QL10 ( .CLK(CLK), .D(N_5), .Q(N_4) );
dff QL11 ( .CLK(CLK), .D(D4), .Q(N_5) );
dff QL12 ( .CLK(CLK), .D(N_1), .Q(N_6) );
dff QL13 ( .CLK(CLK), .D(D3), .Q(N_1) );
dff QL14 ( .CLK(CLK), .D(N_2), .Q(N_7) );
dff QL15 ( .CLK(CLK), .D(D2), .Q(N_2) );
dff QL16 ( .CLK(CLK), .D(D1), .Q(N_3) );

endmodule // ttl396

`endif

`ifdef ttl395q
`else
`define ttl395q
module ttl395q( A , B, C, CLK, CLR, D, LD_SHNN, SER, QA, QB, QC, QD );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input A, B, C, D, LD_SHNN;
output QA, QB, QC, QD;
input SER;
wire N_1;
wire N_2;
wire N_3;
wire N_4;

dffc QL1 ( .CLK(CLK), .CLR(CLR), .D(N_1), .Q(QD) );
dffc QL2 ( .CLK(CLK), .CLR(CLR), .D(N_2), .Q(QC) );
dffc QL3 ( .CLK(CLK), .CLR(CLR), .D(N_3), .Q(QB) );
dffc QL4 ( .CLK(CLK), .CLR(CLR), .D(N_4), .Q(QA) );
mux2x0 QL5 ( .A(QC), .B(D), .Q(N_1), .S(LD_SHNN) );
mux2x0 QL6 ( .A(QB), .B(C), .Q(N_2), .S(LD_SHNN) );
mux2x0 QL7 ( .A(QA), .B(B), .Q(N_3), .S(LD_SHNN) );
mux2x0 QL8 ( .A(SER), .B(A), .Q(N_4), .S(LD_SHNN) );

endmodule // ttl395q

`endif

`ifdef ttl376q
`else
`define ttl376q
module ttl376q( CLK , CLR, J1, J2, J3, J4, KNN1, KNN2, KNN3, KNN4, Q1, Q2, Q3, Q4 );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input J1, J2, J3, J4, KNN1, KNN2, KNN3, KNN4;
output Q1, Q2, Q3, Q4;

jknn_ff QL1 ( .CLK(CLK), .CLR(CLR), .J(J4), .KNN(KNN4), .Q(Q4) );
jknn_ff QL2 ( .CLK(CLK), .CLR(CLR), .J(J3), .KNN(KNN3), .Q(Q3) );
jknn_ff QL3 ( .CLK(CLK), .CLR(CLR), .J(J2), .KNN(KNN2), .Q(Q2) );
jknn_ff QL4 ( .CLK(CLK), .CLR(CLR), .J(J1), .KNN(KNN1), .Q(Q1) );

endmodule // ttl376q

`endif

`ifdef ttl375
`else
`define ttl375
module ttl375( C1_C2 , C3_C4, D1, D2, D3, D4, Q1, Q2, Q3, Q4, QNN1, QNN2, QNN3,
               QNN4 );
input C1_C2, C3_C4, D1, D2, D3, D4;
output Q1, Q2, Q3, Q4, QNN1, QNN2, QNN3, QNN4;

dladinv QL1 ( .DATA(D4), .G(C3_C4), .Q(Q4), .QNN(QNN4) );
dladinv QL2 ( .DATA(D3), .G(C3_C4), .Q(Q3), .QNN(QNN3) );
dladinv QL3 ( .DATA(D2), .G(C1_C2), .Q(Q2), .QNN(QNN2) );
dladinv QL4 ( .DATA(D1), .G(C1_C2), .Q(Q1), .QNN(QNN1) );

endmodule // ttl375

`endif

`ifdef ttl374q
`else
`define ttl374q
module ttl374q( CLK , D1, D2, D3, D4, D5, D6, D7, D8, Q1, Q2, Q3, Q4, Q5, Q6, Q7,
                Q8 );
input CLK /* synthesis syn_isclock=1 */;
input D1, D2, D3, D4, D5, D6, D7, D8;
output Q1, Q2, Q3, Q4, Q5, Q6, Q7, Q8;

dff QL1 ( .CLK(CLK), .D(D8), .Q(Q8) );
dff QL2 ( .CLK(CLK), .D(D7), .Q(Q7) );
dff QL3 ( .CLK(CLK), .D(D6), .Q(Q6) );
dff QL4 ( .CLK(CLK), .D(D5), .Q(Q5) );
dff QL5 ( .CLK(CLK), .D(D4), .Q(Q4) );
dff QL6 ( .CLK(CLK), .D(D3), .Q(Q3) );
dff QL7 ( .CLK(CLK), .D(D2), .Q(Q2) );
dff QL8 ( .CLK(CLK), .D(D1), .Q(Q1) );

endmodule // ttl374q

`endif

`ifdef ttl373q
`else
`define ttl373q
module ttl373q( C , D1, D2, D3, D4, D5, D6, D7, D8, Q1, Q2, Q3, Q4, Q5, Q6, Q7,
                Q8 );
input C, D1, D2, D3, D4, D5, D6, D7, D8;
output Q1, Q2, Q3, Q4, Q5, Q6, Q7, Q8;

dlad QL1 ( .D1(D1), .D2(D2), .G(C), .Q1(Q1), .Q2(Q2) );
dlad QL2 ( .D1(D7), .D2(D8), .G(C), .Q1(Q7), .Q2(Q8) );
dlad QL3 ( .D1(D5), .D2(D6), .G(C), .Q1(Q5), .Q2(Q6) );
dlad QL4 ( .D1(D3), .D2(D4), .G(C), .Q1(Q3), .Q2(Q4) );

endmodule // ttl373q

`endif

`ifdef ttl368
`else
`define ttl368
module ttl368( A1_1 , A1_2, A1_3, A1_4, A2_1, A2_2, GNN1, GNN2, Y1_1, Y1_2, Y1_3,
               Y1_4, Y2_1, Y2_2 );
input A1_1, A1_2, A1_3, A1_4, A2_1, A2_2, GNN1, GNN2;
output Y1_1, Y1_2, Y1_3, Y1_4, Y2_1, Y2_2;
wire N_1;
wire N_2;

inv QL1 ( .A(GNN2), .Q(N_1) );
inv QL2 ( .A(GNN1), .Q(N_2) );
triipad QL3 ( .A(A2_2), .EN(N_1), .P(Y2_2) );
triipad QL4 ( .A(A2_1), .EN(N_1), .P(Y2_1) );
triipad QL5 ( .A(A1_4), .EN(N_2), .P(Y1_4) );
triipad QL6 ( .A(A1_3), .EN(N_2), .P(Y1_3) );
triipad QL7 ( .A(A1_2), .EN(N_2), .P(Y1_2) );
triipad QL8 ( .A(A1_1), .EN(N_2), .P(Y1_1) );

endmodule // ttl368

`endif

`ifdef ttl367
`else
`define ttl367
module ttl367( A1_1 , A1_2, A1_3, A1_4, A2_1, A2_2, GNN1, GNN2, Y1_1, Y1_2, Y1_3,
               Y1_4, Y2_1, Y2_2 );
input A1_1, A1_2, A1_3, A1_4, A2_1, A2_2, GNN1, GNN2;
output Y1_1, Y1_2, Y1_3, Y1_4, Y2_1, Y2_2;
wire N_1;
wire N_2;

inv QL1 ( .A(GNN2), .Q(N_1) );
inv QL2 ( .A(GNN1), .Q(N_2) );
tripad QL3 ( .A(A1_1), .EN(N_2), .P(Y1_1) );
tripad QL4 ( .A(A1_2), .EN(N_2), .P(Y1_2) );
tripad QL5 ( .A(A1_3), .EN(N_2), .P(Y1_3) );
tripad QL6 ( .A(A1_4), .EN(N_2), .P(Y1_4) );
tripad QL7 ( .A(A2_1), .EN(N_1), .P(Y2_1) );
tripad QL8 ( .A(A2_2), .EN(N_1), .P(Y2_2) );

endmodule // ttl367

`endif

`ifdef ttl366
`else
`define ttl366
module ttl366( A1 , A2, A3, A4, A5, A6, G1NN, G2NN, Y1, Y2, Y3, Y4, Y5, Y6 );
input A1, A2, A3, A4, A5, A6, G1NN, G2NN;
output Y1, Y2, Y3, Y4, Y5, Y6;
wire N_1;

triipad QL1 ( .A(A6), .EN(N_1), .P(Y6) );
triipad QL2 ( .A(A5), .EN(N_1), .P(Y5) );
triipad QL3 ( .A(A4), .EN(N_1), .P(Y4) );
triipad QL4 ( .A(A3), .EN(N_1), .P(Y3) );
triipad QL5 ( .A(A2), .EN(N_1), .P(Y2) );
triipad QL6 ( .A(A1), .EN(N_1), .P(Y1) );
and2i2 QL7 ( .A(G1NN), .B(G2NN), .Q(N_1) );

endmodule // ttl366

`endif

`ifdef ttl365
`else
`define ttl365
module ttl365( A1 , A2, A3, A4, A5, A6, G1NN, G2NN, Y1, Y2, Y3, Y4, Y5, Y6 );
input A1, A2, A3, A4, A5, A6, G1NN, G2NN;
output Y1, Y2, Y3, Y4, Y5, Y6;
wire N_1;

and2i2 QL1 ( .A(G1NN), .B(G2NN), .Q(N_1) );
tripad QL2 ( .A(A6), .EN(N_1), .P(Y6) );
tripad QL3 ( .A(A5), .EN(N_1), .P(Y5) );
tripad QL4 ( .A(A2), .EN(N_1), .P(Y2) );
tripad QL5 ( .A(A4), .EN(N_1), .P(Y4) );
tripad QL6 ( .A(A3), .EN(N_1), .P(Y3) );
tripad QL7 ( .A(A1), .EN(N_1), .P(Y1) );

endmodule // ttl365

`endif

`ifdef ttl295q
`else
`define ttl295q
module ttl295q( A , B, C, CLK, D, LD_SHNN, SER, QA, QB, QC, QD );
input CLK /* synthesis syn_isclock=1 */;
input A, B, C, D, LD_SHNN;
output QA, QB, QC, QD;
input SER;
wire N_1;
wire N_2;
wire N_3;
wire N_4;

mux2x0 QL1 ( .A(QC), .B(D), .Q(N_1), .S(LD_SHNN) );
mux2x0 QL2 ( .A(QB), .B(C), .Q(N_2), .S(LD_SHNN) );
mux2x0 QL3 ( .A(QA), .B(B), .Q(N_3), .S(LD_SHNN) );
mux2x0 QL4 ( .A(SER), .B(A), .Q(N_4), .S(LD_SHNN) );
dff QL5 ( .CLK(CLK), .D(N_3), .Q(QB) );
dff QL6 ( .CLK(CLK), .D(N_4), .Q(QA) );
dff QL7 ( .CLK(CLK), .D(N_1), .Q(QD) );
dff QL8 ( .CLK(CLK), .D(N_2), .Q(QC) );

endmodule // ttl295q

`endif

`ifdef ttl279
`else
`define ttl279
module ttl279( RNN1 , RNN2, RNN3, RNN4, S1NN1, S1NN3, S2NN1, S2NN3, SNN2, SNN4, Q1,
               Q2, Q3, Q4 );
output Q1, Q2, Q3, Q4;
input RNN1, RNN2, RNN3, RNN4, S1NN1, S1NN3, S2NN1, S2NN3, SNN2, SNN4;

s_r_ltch I_1 ( .Q(Q4), .R(RNN4), .S1(SNN4), .S2(SNN4) );
s_r_ltch I_2 ( .Q(Q3), .R(RNN3), .S1(S1NN3), .S2(S2NN3) );
s_r_ltch I_3 ( .Q(Q2), .R(RNN2), .S1(SNN2), .S2(SNN2) );
s_r_ltch I_4 ( .Q(Q1), .R(RNN1), .S1(S1NN1), .S2(S2NN1) );

endmodule // ttl279

`endif

`ifdef ttl278
`else
`define ttl278
module ttl278( D1 , D2, D3, D4, G, P0, P1, Y1, Y2, Y3, Y4 );
input D1, D2, D3, D4, G, P0;
output P1, Y1, Y2, Y3, Y4;
wire N_1;
wire N_2;
wire N_3;
wire N_4;

ttl77 QL1 ( .C1C2(G), .C3C4(G), .D1(D1), .D2(D2), .D3(D3), .D4(D4), .Q1(N_4),
         .Q2(N_3), .Q3(N_2), .Q4(N_1) );
or5i0 QL2 ( .A(P0), .B(N_4), .C(N_3), .D(N_2), .E(N_1), .Q(P1) );
nor5i1 QL3 ( .A(P0), .B(N_4), .C(N_3), .D(N_2), .E(N_1), .Q(Y4) );
nor4i1 QL4 ( .A(P0), .B(N_4), .C(N_3), .D(N_2), .Q(Y3) );
nor3i1 QL5 ( .A(P0), .B(N_4), .C(N_3), .Q(Y2) );
nor2i1 QL6 ( .A(P0), .B(N_4), .Q(Y1) );

endmodule // ttl278

`endif

`ifdef ttl273q
`else
`define ttl273q
module ttl273q( CLEAR , CLK, D1, D2, D3, D4, D5, D6, D7, D8, Q1, Q2, Q3, Q4, Q5, Q6,
                Q7, Q8 );
input CLK /* synthesis syn_isclock=1 */;
input CLEAR /* synthesis syn_isclock=1 */;
input D1, D2, D3, D4, D5, D6, D7, D8;
output Q1, Q2, Q3, Q4, Q5, Q6, Q7, Q8;

dffc QL1 ( .CLK(CLK), .CLR(CLEAR), .D(D8), .Q(Q8) );
dffc QL2 ( .CLK(CLK), .CLR(CLEAR), .D(D7), .Q(Q7) );
dffc QL3 ( .CLK(CLK), .CLR(CLEAR), .D(D6), .Q(Q6) );
dffc QL4 ( .CLK(CLK), .CLR(CLEAR), .D(D5), .Q(Q5) );
dffc QL5 ( .CLK(CLK), .CLR(CLEAR), .D(D4), .Q(Q4) );
dffc QL6 ( .CLK(CLK), .CLR(CLEAR), .D(D3), .Q(Q3) );
dffc QL7 ( .CLK(CLK), .CLR(CLEAR), .D(D2), .Q(Q2) );
dffc QL8 ( .CLK(CLK), .CLR(CLEAR), .D(D1), .Q(Q1) );

endmodule // ttl273q

`endif

`ifdef ttl27
`else
`define ttl27
module ttl27( A1 , A2, A3, B1, B2, B3, C1, C2, C3, Y1, Y2, Y3 );
input A1, A2, A3, B1, B2, B3, C1, C2, C3;
output Y1, Y2, Y3;

nor3i0 QL1 ( .A(A1), .B(B1), .C(C1), .Q(Y1) );
nor3i0 QL2 ( .A(A2), .B(B2), .C(C2), .Q(Y2) );
nor3i0 QL3 ( .A(A3), .B(B3), .C(C3), .Q(Y3) );

endmodule // ttl27

`endif

`ifdef ttl268q
`else
`define ttl268q
module ttl268q( C , D1, D2, D3, D4, D5, D6, Q1, Q2, Q3, Q4, Q5, Q6 );
input C, D1, D2, D3, D4, D5, D6;
output Q1, Q2, Q3, Q4, Q5, Q6;

dlad QL1 ( .D1(D5), .D2(D6), .G(C), .Q1(Q5), .Q2(Q6) );
dlad QL2 ( .D1(D3), .D2(D4), .G(C), .Q1(Q3), .Q2(Q4) );
dlad QL3 ( .D1(D1), .D2(D2), .G(C), .Q1(Q1), .Q2(Q2) );

endmodule // ttl268q

`endif

`ifdef ttl259
`else
`define ttl259
module ttl259( CLRNN , DATA, GNN, S0, S1, S2, Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7 );
input CLRNN, DATA, GNN;
output Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7;
input S0, S1, S2;
wire N_1;
supply0 GND;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;

bank259 I_1 ( .CLRNN(CLRNN), .D0(N_8), .D1(N_7), .D2(N_6), .D3(N_5), .D4(N_4),
           .D5(N_3), .D6(N_1), .D7(N_2), .DATA(DATA), .GNN(GNN), .Q0(Q0),
           .Q1(Q1), .Q2(Q2), .Q3(Q3), .Q4(Q4), .Q5(Q5), .Q6(Q6), .Q7(Q7) );
ttl138q QL1 ( .A(S0), .B(S1), .C(S2), .EN(GND), .Y0(N_8), .Y1(N_7), .Y2(N_6),
           .Y3(N_5), .Y4(N_4), .Y5(N_3), .Y6(N_1), .Y7(N_2) );

endmodule // ttl259

`endif

`ifdef ttl244q
`else
`define ttl244q
module ttl244q( A1_1 , A1_2, A1_3, A1_4, A2_1, A2_2, A2_3, A2_4, G1, G2, Y1_1,
                Y1_2, Y1_3, Y1_4, Y2_1, Y2_2, Y2_3, Y2_4 );
input A1_1, A1_2, A1_3, A1_4, A2_1, A2_2, A2_3, A2_4, G1, G2;
output Y1_1, Y1_2, Y1_3, Y1_4, Y2_1, Y2_2, Y2_3, Y2_4;

tripad QL1 ( .A(A2_4), .EN(G2), .P(Y2_4) );
tripad QL2 ( .A(A2_3), .EN(G2), .P(Y2_3) );
tripad QL3 ( .A(A2_2), .EN(G2), .P(Y2_2) );
tripad QL4 ( .A(A2_1), .EN(G2), .P(Y2_1) );
tripad QL5 ( .A(A1_4), .EN(G1), .P(Y1_4) );
tripad QL6 ( .A(A1_3), .EN(G1), .P(Y1_3) );
tripad QL7 ( .A(A1_2), .EN(G1), .P(Y1_2) );
tripad QL8 ( .A(A1_1), .EN(G1), .P(Y1_1) );

endmodule // ttl244q

`endif

`ifdef ttl240q
`else
`define ttl240q
module ttl240q( A1_1 , A1_2, A1_3, A1_4, A2_1, A2_2, A2_3, A2_4, G1, G2, Y1, Y2 );
input A1_1, A1_2, A1_3, A1_4, A2_1, A2_2, A2_3, A2_4, G1, G2;
 output [4:1] Y1;
 output [4:1] Y2;

triipad QL1 ( .A(A1_4), .EN(G1), .P(Y1[4]) );
triipad QL2 ( .A(A1_3), .EN(G1), .P(Y1[3]) );
triipad QL3 ( .A(A1_2), .EN(G1), .P(Y1[2]) );
triipad QL4 ( .A(A1_1), .EN(G1), .P(Y1[1]) );
triipad QL5 ( .A(A2_4), .EN(G2), .P(Y2[4]) );
triipad QL6 ( .A(A2_3), .EN(G2), .P(Y2[3]) );
triipad QL7 ( .A(A2_2), .EN(G2), .P(Y2[2]) );
triipad QL8 ( .A(A2_1), .EN(G2), .P(Y2[1]) );

endmodule // ttl240q

`endif

`ifdef ttl21
`else
`define ttl21
module ttl21( A1 , A2, B1, B2, C1, C2, D1, D2, Y1, Y2 );
input A1, A2, B1, B2, C1, C2, D1, D2;
output Y1, Y2;

and4i0 QL1 ( .A(A2), .B(B2), .C(C2), .D(D2), .Q(Y2) );
and4i0 QL2 ( .A(A1), .B(B1), .C(C1), .D(D1), .Q(Y1) );

endmodule // ttl21

`endif

`ifdef ttl194q
`else
`define ttl194q
module ttl194q( A , B, C, CLK, CLR, D, S0, S1, SHFTINL, SHFTINR, QA, QB, QC, QD );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input A, B, C, D;
output QA, QB, QC, QD;
input S0, S1, SHFTINL, SHFTINR;
wire N_1;
wire N_2;
wire N_3;
wire N_4;

dffc QL1 ( .CLK(CLK), .CLR(CLR), .D(N_1), .Q(QA) );
dffc QL2 ( .CLK(CLK), .CLR(CLR), .D(N_4), .Q(QB) );
dffc QL3 ( .CLK(CLK), .CLR(CLR), .D(N_3), .Q(QC) );
dffc QL4 ( .CLK(CLK), .CLR(CLR), .D(N_2), .Q(QD) );
mux4x0 QL5 ( .A(QA), .B(SHFTINR), .C(QB), .D(A), .Q(N_1), .S0(S0), .S1(S1) );
mux4x0 QL6 ( .A(QB), .B(QA), .C(QC), .D(B), .Q(N_4), .S0(S0), .S1(S1) );
mux4x0 QL7 ( .A(QC), .B(QB), .C(QD), .D(C), .Q(N_3), .S0(S0), .S1(S1) );
mux4x0 QL8 ( .A(QD), .B(QC), .C(SHFTINL), .D(D), .Q(N_2), .S0(S0), .S1(S1) );

endmodule // ttl194q

`endif

`ifdef ttl180
`else
`define ttl180
module ttl180( A , B, C, D, E, EVENIN, F, G, H, ODDIN, EVENOUT, ODDOUT );
input A, B, C, D, E, EVENIN;
output EVENOUT;
input F, G, H, ODDIN;
output ODDOUT;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;

and2i2 QL1 ( .A(N_2), .B(N_1), .Q(ODDOUT) );
and2i2 QL2 ( .A(N_4), .B(N_3), .Q(EVENOUT) );
and2i1 QL3 ( .A(ODDIN), .B(N_5), .Q(N_1) );
and2i1 QL4 ( .A(EVENIN), .B(N_5), .Q(N_3) );
and2i0 QL5 ( .A(N_5), .B(ODDIN), .Q(N_4) );
and2i0 QL6 ( .A(EVENIN), .B(N_5), .Q(N_2) );
xnor2i0 QL7 ( .A(N_6), .B(N_7), .Q(N_5) );
xor3i0 QL8 ( .A(D), .B(E), .C(F), .Q(N_8) );
xor3i0 QL9 ( .A(N_8), .B(G), .C(H), .Q(N_7) );
xor3i0 QL10 ( .A(A), .B(B), .C(C), .Q(N_6) );

endmodule // ttl180

`endif

`ifdef ttl174q
`else
`define ttl174q
module ttl174q( CLK , CLR, D1, D2, D3, D4, D5, D6, Q1, Q2, Q3, Q4, Q5, Q6 );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input D1, D2, D3, D4, D5, D6;
output Q1, Q2, Q3, Q4, Q5, Q6;

dffc QL1 ( .CLK(CLK), .CLR(CLR), .D(D6), .Q(Q6) );
dffc QL2 ( .CLK(CLK), .CLR(CLR), .D(D5), .Q(Q5) );
dffc QL3 ( .CLK(CLK), .CLR(CLR), .D(D4), .Q(Q4) );
dffc QL4 ( .CLK(CLK), .CLR(CLR), .D(D1), .Q(Q1) );
dffc QL5 ( .CLK(CLK), .CLR(CLR), .D(D3), .Q(Q3) );
dffc QL6 ( .CLK(CLK), .CLR(CLR), .D(D2), .Q(Q2) );

endmodule // ttl174q

`endif

`ifdef ttl171q
`else
`define ttl171q
module ttl171q( CLK , CLR, D1, D2, D3, D4, Q1, Q2, Q3, Q4 );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input D1, D2, D3, D4;
output Q1, Q2, Q3, Q4;

dffc QL1 ( .CLK(CLK), .CLR(CLR), .D(D1), .Q(Q1) );
dffc QL2 ( .CLK(CLK), .CLR(CLR), .D(D4), .Q(Q4) );
dffc QL3 ( .CLK(CLK), .CLR(CLR), .D(D3), .Q(Q3) );
dffc QL4 ( .CLK(CLK), .CLR(CLR), .D(D2), .Q(Q2) );

endmodule // ttl171q

`endif

`ifdef ttl169
`else
`define ttl169
module ttl169( CLK , DA, DB, DC, DD, ENPNN, ENTNN, LDNN, UPDWN, QA, QB, QC, QD,
               RCO );
input CLK /* synthesis syn_isclock=1 */;
input DA, DB, DC, DD, ENPNN, ENTNN, LDNN;
output QA, QB, QC, QD, RCO;
input UPDWN;
wire N_1;
wire N_2;
supply0 GND;
wire N_3;
wire N_4;
wire N_5;
wire N_6;

a169 I_1 ( .A(N_4), .ANN(N_5), .OUTB(N_3), .QA(QA), .QB(QB), .UPDWN(UPDWN) );
b169 I_2 ( .A(N_4), .ANN(N_5), .OUTC(N_6), .QC(QC) );
rco169 I_3 ( .A(N_4), .ANN(N_5), .ENT(ENTNN), .QC(QC), .QD(QD), .RCO(RCO) );
reg169 I_4 ( .CLK(CLK), .D_IN(DD), .DATA(N_6), .EN(N_2), .FDBK(QD), .LDNN(LDNN),
          .Q(QD) );
reg169 I_5 ( .CLK(CLK), .D_IN(DC), .DATA(N_3), .EN(N_2), .FDBK(QC), .LDNN(LDNN),
          .Q(QC) );
reg169 I_6 ( .CLK(CLK), .D_IN(DB), .DATA(N_1), .EN(N_2), .FDBK(QB), .LDNN(LDNN),
          .Q(QB) );
reg169 I_7 ( .CLK(CLK), .D_IN(DA), .DATA(GND), .EN(N_2), .FDBK(QA), .LDNN(LDNN),
          .Q(QA) );
mux2x2 QL4 ( .A(QA), .B(QA), .Q(N_1), .S(UPDWN) );
and2i2 QL5 ( .A(ENTNN), .B(ENPNN), .Q(N_2) );

endmodule // ttl169

`endif

`ifdef ttl166q
`else
`define ttl166q
module ttl166q( A , B, C, CLK, CLR, D, E, F, G, H, SER_IN, SH_LDNN, QH );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input A, B, C, D, E, F, G, H;
output QH;
input SER_IN, SH_LDNN;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;
wire N_15;

dffc QL1 ( .CLK(CLK), .CLR(CLR), .D(N_5), .Q(QH) );
dffc QL2 ( .CLK(CLK), .CLR(CLR), .D(N_6), .Q(N_3) );
dffc QL3 ( .CLK(CLK), .CLR(CLR), .D(N_7), .Q(N_4) );
dffc QL4 ( .CLK(CLK), .CLR(CLR), .D(N_8), .Q(N_2) );
dffc QL5 ( .CLK(CLK), .CLR(CLR), .D(N_9), .Q(N_1) );
dffc QL6 ( .CLK(CLK), .CLR(CLR), .D(N_13), .Q(N_10) );
dffc QL7 ( .CLK(CLK), .CLR(CLR), .D(N_14), .Q(N_11) );
dffc QL8 ( .CLK(CLK), .CLR(CLR), .D(N_15), .Q(N_12) );
mux2x0 QL9 ( .A(H), .B(N_3), .Q(N_5), .S(SH_LDNN) );
mux2x0 QL10 ( .A(G), .B(N_4), .Q(N_6), .S(SH_LDNN) );
mux2x0 QL11 ( .A(F), .B(N_2), .Q(N_7), .S(SH_LDNN) );
mux2x0 QL12 ( .A(E), .B(N_1), .Q(N_8), .S(SH_LDNN) );
mux2x0 QL13 ( .A(D), .B(N_10), .Q(N_9), .S(SH_LDNN) );
mux2x0 QL14 ( .A(C), .B(N_11), .Q(N_13), .S(SH_LDNN) );
mux2x0 QL15 ( .A(B), .B(N_12), .Q(N_14), .S(SH_LDNN) );
mux2x0 QL16 ( .A(A), .B(SER_IN), .Q(N_15), .S(SH_LDNN) );

endmodule // ttl166q

`endif

`ifdef ttl164q
`else
`define ttl164q
module ttl164q( A , B, CLK, CLR, QA, QB, QC, QD, QE, QF, QG, QH );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input A, B;
output QA, QB, QC, QD, QE, QF, QG, QH;
wire N_1;

and2i0 QL1 ( .A(A), .B(B), .Q(N_1) );
dffc QL2 ( .CLK(CLK), .CLR(CLR), .D(QG), .Q(QH) );
dffc QL3 ( .CLK(CLK), .CLR(CLR), .D(QF), .Q(QG) );
dffc QL4 ( .CLK(CLK), .CLR(CLR), .D(QE), .Q(QF) );
dffc QL5 ( .CLK(CLK), .CLR(CLR), .D(QD), .Q(QE) );
dffc QL6 ( .CLK(CLK), .CLR(CLR), .D(QC), .Q(QD) );
dffc QL7 ( .CLK(CLK), .CLR(CLR), .D(QB), .Q(QC) );
dffc QL8 ( .CLK(CLK), .CLR(CLR), .D(QA), .Q(QB) );
dffc QL9 ( .CLK(CLK), .CLR(CLR), .D(N_1), .Q(QA) );

endmodule // ttl164q

`endif

`ifdef ttl163
`else
`define ttl163
module ttl163( CLK , CLR, D, ENP, ENT, LOAD, Q, RCO );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [3:0] D;
input ENP, ENT, LOAD;
 output [3:0] Q;
output RCO;
supply1 VCC;

uplsbit QL1 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(VCC) );
uplsbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
uplsbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[1]), .Q0(Q[0]), .Q1(VCC), .Q2(VCC) );
uplsbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[0]), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
nand5i1 QL5 ( .A(Q[0]), .B(Q[1]), .C(Q[2]), .D(Q[3]), .E(ENT), .Q(RCO) );

endmodule // ttl163

`endif

`ifdef ttl161
`else
`define ttl161
module ttl161( CLK , CLR, D, ENP, ENT, LOAD, Q, RCO );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [3:0] D;
input ENP, ENT, LOAD;
 output [3:0] Q;
output RCO;
supply1 VCC;

uplabit QL1 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
uplabit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(VCC) );
uplabit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[1]), .Q0(Q[0]), .Q1(VCC), .Q2(VCC) );
uplabit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[0]), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
nand5i1 QL5 ( .A(Q[0]), .B(Q[1]), .C(Q[2]), .D(Q[3]), .E(ENT), .Q(RCO) );

endmodule // ttl161

`endif

`ifdef ttl157
`else
`define ttl157
module ttl157( A1 , A2, A3, A4, B1, B2, B3, B4, SEL, STRBNN, Y1, Y2, Y3, Y4 );
input A1, A2, A3, A4, B1, B2, B3, B4, SEL, STRBNN;
output Y1, Y2, Y3, Y4;

muxde2x0 QL1 ( .A1(A3), .A2(A4), .B1(B3), .B2(B4), .GNN(STRBNN), .SEL(SEL), .Y1(Y3),
            .Y2(Y4) );
muxde2x0 QL2 ( .A1(A1), .A2(A2), .B1(B1), .B2(B2), .GNN(STRBNN), .SEL(SEL), .Y1(Y1),
            .Y2(Y2) );

endmodule // ttl157

`endif

`ifdef ttl154q
`else
`define ttl154q
module ttl154q( A , B, C, D, G1NN, G2NN, Q0, Q1, Q10, Q11, Q12, Q13, Q14, Q15,
                Q2, Q3, Q4, Q5, Q6, Q7, Q8, Q9 );
input A, B, C, D, G1NN, G2NN;
output Q0, Q1, Q10, Q11, Q12, Q13, Q14, Q15, Q2, Q3, Q4, Q5, Q6, Q7, Q8, Q9;

and6i2 QL1 ( .A(A), .B(B), .C(C), .D(D), .E(G1NN), .F(G2NN), .Q(Q15) );
and6i3 QL2 ( .A(B), .B(C), .C(D), .D(A), .E(G1NN), .F(G2NN), .Q(Q14) );
and6i3 QL3 ( .A(A), .B(C), .C(D), .D(B), .E(G1NN), .F(G2NN), .Q(Q13) );
and6i3 QL4 ( .A(A), .B(B), .C(D), .D(C), .E(G1NN), .F(G2NN), .Q(Q11) );
and6i3 QL5 ( .A(A), .B(B), .C(C), .D(D), .E(G1NN), .F(G2NN), .Q(Q7) );
and6i4 QL6 ( .A(C), .B(D), .C(A), .D(B), .E(G1NN), .F(G2NN), .Q(Q12) );
and6i4 QL7 ( .A(B), .B(D), .C(A), .D(C), .E(G1NN), .F(G2NN), .Q(Q10) );
and6i4 QL8 ( .A(A), .B(D), .C(B), .D(C), .E(G1NN), .F(G2NN), .Q(Q9) );
and6i4 QL9 ( .A(B), .B(C), .C(A), .D(D), .E(G1NN), .F(G2NN), .Q(Q6) );
and6i4 QL10 ( .A(A), .B(C), .C(B), .D(D), .E(G1NN), .F(G2NN), .Q(Q5) );
and6i4 QL11 ( .A(A), .B(B), .C(C), .D(D), .E(G1NN), .F(G2NN), .Q(Q3) );
and6i5 QL12 ( .A(D), .B(A), .C(B), .D(C), .E(G1NN), .F(G2NN), .Q(Q8) );
and6i5 QL13 ( .A(C), .B(A), .C(B), .D(D), .E(G1NN), .F(G2NN), .Q(Q4) );
and6i5 QL14 ( .A(B), .B(A), .C(C), .D(D), .E(G1NN), .F(G2NN), .Q(Q2) );
and6i5 QL15 ( .A(A), .B(B), .C(C), .D(D), .E(G1NN), .F(G2NN), .Q(Q1) );
and6i6 QL16 ( .A(A), .B(B), .C(C), .D(D), .E(G1NN), .F(G2NN), .Q(Q0) );

endmodule // ttl154q

`endif

`ifdef ttl153
`else
`define ttl153
module ttl153( C1_0 , C1_1, C1_2, C1_3, C2_0, C2_1, C2_2, C2_3, GNN1, GNN2, S0, S1,
               Y1, Y2 );
input C1_0, C1_1, C1_2, C1_3, C2_0, C2_1, C2_2, C2_3, GNN1, GNN2, S0, S1;
output Y1, Y2;

mux4x0e QL1 ( .A(C2_0), .B(C2_1), .C(C2_2), .D(C2_3), .GNN(GNN2), .Q(Y2), .S0(S0),
           .S1(S1) );
mux4x0e QL2 ( .A(C1_0), .B(C1_1), .C(C1_2), .D(C1_3), .GNN(GNN1), .Q(Y1), .S0(S0),
           .S1(S1) );

endmodule // ttl153

`endif

`ifdef ttl152
`else
`define ttl152
module ttl152( A , B, C, D0, D1, D2, D3, D4, D5, D6, D7, W );
input A, B, C, D0, D1, D2, D3, D4, D5, D6, D7;
output W;
wire N_1;
wire N_2;

mux4x0 QL1 ( .A(D0), .B(D1), .C(D2), .D(D3), .Q(N_1), .S0(A), .S1(B) );
mux4x0 QL2 ( .A(D4), .B(D5), .C(D6), .D(D7), .Q(N_2), .S0(A), .S1(B) );
mux2x0 QL3 ( .A(N_1), .B(N_2), .Q(W), .S(C) );

endmodule // ttl152

`endif

`ifdef ttl150
`else
`define ttl150
module ttl150( A , B, C, D, E0, E1, E10, E11, E12, E13, E14, E15, E2, E3, E4,
               E5, E6, E7, E8, E9, STRBNN, W );
input A, B, C, D, E0, E1, E10, E11, E12, E13, E14, E15, E2, E3, E4, E5, E6,
E7, E8, E9, STRBNN;
output W;
supply1 VCC;
supply0 GND;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;
wire N_15;
wire N_16;
wire N_17;
wire N_18;
wire N_19;
wire N_20;
wire N_21;

and14i7 QL1 ( .A(N_11), .B(N_10), .C(N_9), .D(N_1), .E(N_2), .F(VCC), .G(VCC),
           .H(GND), .I(N_7), .J(N_8), .K(N_3), .L(N_4), .M(N_5), .N(N_6), .Q(W) );
nor2i0 QL2 ( .A(N_13), .B(N_12), .Q(N_2) );
nor2i0 QL3 ( .A(N_15), .B(N_14), .Q(N_1) );
nor2i0 QL4 ( .A(N_17), .B(N_16), .Q(N_9) );
nor2i0 QL5 ( .A(N_19), .B(N_18), .Q(N_10) );
nor2i0 QL6 ( .A(N_21), .B(N_20), .Q(N_11) );
and6i1 QL7 ( .A(E15), .B(A), .C(B), .D(C), .E(D), .F(STRBNN), .Q(N_6) );
and6i2 QL8 ( .A(E14), .B(B), .C(C), .D(D), .E(A), .F(STRBNN), .Q(N_5) );
and6i2 QL9 ( .A(E13), .B(A), .C(C), .D(D), .E(B), .F(STRBNN), .Q(N_4) );
and6i2 QL10 ( .A(E11), .B(A), .C(B), .D(D), .E(C), .F(STRBNN), .Q(N_12) );
and6i2 QL11 ( .A(E7), .B(A), .C(B), .D(C), .E(D), .F(STRBNN), .Q(N_16) );
and6i3 QL12 ( .A(E12), .B(C), .C(D), .D(A), .E(B), .F(STRBNN), .Q(N_3) );
and6i3 QL13 ( .A(E10), .B(B), .C(D), .D(A), .E(C), .F(STRBNN), .Q(N_13) );
and6i3 QL14 ( .A(E9), .B(A), .C(D), .D(B), .E(C), .F(STRBNN), .Q(N_14) );
and6i3 QL15 ( .A(E6), .B(B), .C(C), .D(A), .E(D), .F(STRBNN), .Q(N_17) );
and6i3 QL16 ( .A(E5), .B(A), .C(C), .D(B), .E(D), .F(STRBNN), .Q(N_18) );
and6i3 QL17 ( .A(E3), .B(A), .C(B), .D(C), .E(D), .F(STRBNN), .Q(N_20) );
and6i4 QL18 ( .A(E8), .B(D), .C(A), .D(B), .E(C), .F(STRBNN), .Q(N_15) );
and6i4 QL19 ( .A(E4), .B(C), .C(A), .D(B), .E(D), .F(STRBNN), .Q(N_19) );
and6i4 QL20 ( .A(E2), .B(B), .C(A), .D(C), .E(D), .F(STRBNN), .Q(N_21) );
and6i4 QL21 ( .A(E1), .B(A), .C(B), .D(C), .E(D), .F(STRBNN), .Q(N_8) );
and6i5 QL22 ( .A(E0), .B(A), .C(B), .D(C), .E(D), .F(STRBNN), .Q(N_7) );

endmodule // ttl150

`endif

`ifdef ttl148
`else
`define ttl148
module ttl148( EI , P0, P1, P2, P3, P4, P5, P6, P7, A0, A1, A2, EO, GS );
output A0, A1, A2;
input EI;
output EO, GS;
input P0, P1, P2, P3, P4, P5, P6, P7;
wire N_1;

t148a2 I_2 ( .A2(A2), .EI(EI), .P4(P4), .P5(P5), .P6(P6), .P7(P7) );
t148a1 I_3 ( .A1(A1), .EI(EI), .P2(P3), .P3(P2), .P4(P4), .P5(P5), .P6(P6), .P7(P7) );
t148ao I_1 ( .A0(A0), .EI(EI), .P1(P1), .P2(P2), .P3(P3), .P4(P4), .P5(P5), .P6(P6),
          .P7(P7) );
nand4i1 QL1 ( .A(N_1), .B(P6), .C(P7), .D(EI), .Q(EO) );
and6i0 QL2 ( .A(P1), .B(P2), .C(P3), .D(P4), .E(P5), .F(P0), .Q(N_1) );
nand2i1 QL3 ( .A(EO), .B(EI), .Q(GS) );

endmodule // ttl148

`endif

`ifdef ttl145q
`else
`define ttl145q
module ttl145q( INA , INB, INC, IND, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5, OUT6,
                OUT7, OUT8, OUT9 );
input INA, INB, INC, IND;
output OUT0, OUT1, OUT2, OUT3, OUT4, OUT5, OUT6, OUT7, OUT8, OUT9;

and4i1 QL1 ( .A(INA), .B(INB), .C(INC), .D(IND), .Q(OUT7) );
and4i2 QL2 ( .A(IND), .B(INA), .C(INB), .D(INC), .Q(OUT9) );
and4i2 QL3 ( .A(INB), .B(INC), .C(INA), .D(IND), .Q(OUT6) );
and4i2 QL4 ( .A(INA), .B(INC), .C(INB), .D(IND), .Q(OUT5) );
and4i2 QL5 ( .A(INA), .B(INB), .C(INC), .D(IND), .Q(OUT3) );
and4i3 QL6 ( .A(IND), .B(INA), .C(INB), .D(INC), .Q(OUT8) );
and4i3 QL7 ( .A(INA), .B(INB), .C(INC), .D(IND), .Q(OUT1) );
and4i3 QL8 ( .A(INC), .B(INA), .C(INB), .D(IND), .Q(OUT4) );
and4i3 QL9 ( .A(INB), .B(INA), .C(INC), .D(IND), .Q(OUT2) );
and4i4 QL10 ( .A(INA), .B(INB), .C(INC), .D(IND), .Q(OUT0) );

endmodule // ttl145q

`endif

`ifdef ttl139q
`else
`define ttl139q
module ttl139q( A1 , A2, B1, B2, GNN1, GNN2, Y1_0, Y1_1, Y1_2, Y1_3, Y2_0, Y2_1,
                Y2_2, Y2_3 );
input A1, A2, B1, B2, GNN1, GNN2;
output Y1_0, Y1_1, Y1_2, Y1_3, Y2_0, Y2_1, Y2_2, Y2_3;

and3i1 QL1 ( .A(A2), .B(B2), .C(GNN2), .Q(Y2_3) );
and3i1 QL2 ( .A(A1), .B(B1), .C(GNN1), .Q(Y1_3) );
and3i2 QL3 ( .A(B2), .B(A2), .C(GNN2), .Q(Y2_2) );
and3i2 QL4 ( .A(A2), .B(B2), .C(GNN2), .Q(Y2_1) );
and3i2 QL5 ( .A(B1), .B(A1), .C(GNN1), .Q(Y1_2) );
and3i2 QL6 ( .A(A1), .B(B1), .C(GNN1), .Q(Y1_1) );
and3i3 QL7 ( .A(A2), .B(B2), .C(GNN2), .Q(Y2_0) );
and3i3 QL8 ( .A(A1), .B(B1), .C(GNN1), .Q(Y1_0) );

endmodule // ttl139q

`endif

`ifdef ttl138q
`else
`define ttl138q
module ttl138q( A , B, C, EN, Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7 );
input A, B, C, EN;
output Y0, Y1, Y2, Y3, Y4, Y5, Y6, Y7;
wire N_1;

t138f3 I_1 ( .A(A), .B(B), .C(C), .EN(EN), .ENOUT(N_1), .Y1(Y1), .Y5(Y5) );
t138f2 I_2 ( .A(A), .B(B), .C(C), .EN(N_1), .Y0(Y0), .Y3(Y3), .Y6(Y6) );
t138f1 I_3 ( .A(A), .B(B), .C(C), .EN(EN), .Y2(Y2), .Y4(Y4), .Y7(Y7) );

endmodule // ttl138q

`endif

`ifdef ttl116
`else
`define ttl116
module ttl116( C1NN1 , C1NN2, C2NN1, C2NN2, CLR1, CLR2, D1_1, D1_2, D1_3, D1_4,
               D2_1, D2_2, D2_3, D2_4, Q1_1, Q1_2, Q1_3, Q1_4, Q2_1, Q2_2,
               Q2_3, Q2_4 );
input CLR1 /* synthesis syn_isclock=1 */;
input CLR2 /* synthesis syn_isclock=1 */;
input C1NN1, C1NN2, C2NN1, C2NN2, D1_1, D1_2, D1_3, D1_4, D2_1,
D2_2, D2_3, D2_4;
output Q1_1, Q1_2, Q1_3, Q1_4, Q2_1, Q2_2, Q2_3, Q2_4;

dladc QL1 ( .C1NN(C1NN2), .C2NN(C2NN2), .CLR(CLR2), .D1(D2_3), .D2(D2_4),
         .Q1(Q2_3), .Q2(Q2_4) );
dladc QL2 ( .C1NN(C1NN2), .C2NN(C2NN2), .CLR(CLR2), .D1(D2_1), .D2(D2_2),
         .Q1(Q2_1), .Q2(Q2_2) );
dladc QL3 ( .C1NN(C1NN1), .C2NN(C2NN1), .CLR(CLR1), .D1(D1_3), .D2(D1_4),
         .Q1(Q1_3), .Q2(Q1_4) );
dladc QL4 ( .C1NN(C1NN1), .C2NN(C2NN1), .CLR(CLR1), .D1(D1_1), .D2(D1_2),
         .Q1(Q1_1), .Q2(Q1_2) );

endmodule // ttl116

`endif

`ifdef ttl11
`else
`define ttl11
module ttl11( A1 , A2, A3, B1, B2, B3, C1, C2, C3, Y1, Y2, Y3 );
input A1, A2, A3, B1, B2, B3, C1, C2, C3;
output Y1, Y2, Y3;

and3i0 QL1 ( .A(A3), .B(B3), .C(C3), .Q(Y3) );
and3i0 QL2 ( .A(A2), .B(B2), .C(C2), .Q(Y2) );
and3i0 QL3 ( .A(A1), .B(B1), .C(C1), .Q(Y1) );

endmodule // ttl11

`endif

`ifdef ttl109q
`else
`define ttl109q
module ttl109q( CLK1 , CLK2, CLR1, CLR2, J1, J2, KNN1, KNN2, PRE1, PRE2, Q1, Q2 );
input CLK1 /* synthesis syn_isclock=1 */;
input CLK2 /* synthesis syn_isclock=1 */;
input CLR1 /* synthesis syn_isclock=1 */;
input CLR2 /* synthesis syn_isclock=1 */;
input PRE1 /* synthesis syn_isclock=1 */;
input PRE2 /* synthesis syn_isclock=1 */;
input J1, J2, KNN1, KNN2;
output Q1, Q2;

jknffpc QL1 ( .CLK(CLK2), .CLR(CLR2), .J(J2), .K(KNN2), .PRE(PRE2), .Q(Q2) );
jknffpc QL2 ( .CLK(CLK1), .CLR(CLR1), .J(J1), .K(KNN1), .PRE(PRE1), .Q(Q1) );

endmodule // ttl109q

`endif

`ifdef ttl107q
`else
`define ttl107q
module ttl107q( CLK1 , CLK2, CLR1, CLR2, J1, J2, K1, K2, Q1, Q2 );
input CLK1 /* synthesis syn_isclock=1 */;
input CLK2 /* synthesis syn_isclock=1 */;
input CLR1 /* synthesis syn_isclock=1 */;
input CLR2 /* synthesis syn_isclock=1 */;
input J1, J2, K1, K2;
output Q1, Q2;
supply0 GND;

jkffpc QL1 ( .CLK(CLK2), .CLR(CLR2), .J(J2), .K(K2), .PRE(GND), .Q(Q2) );
jkffpc QL2 ( .CLK(CLK1), .CLR(CLR1), .J(J1), .K(K1), .PRE(GND), .Q(Q1) );

endmodule // ttl107q

`endif

`ifdef ttl105q
`else
`define ttl105q
module ttl105q( CLK , CLR, J1, J2NN, J3, JK, K1, K2NN, K3, PRE, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input PRE /* synthesis syn_isclock=1 */;
input J1, J2NN, J3, JK, K1, K2NN, K3;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(PRE), .QZ(Q) );
frag_f I_2 ( .F1(K1), .F2(K2NN), .F3(JK), .F4(GND), .F5(K3), .F6(GND), .FZ(N_3) );
frag_m I_1 ( .B1(Q), .B2(GND), .C1(GND), .C2(VCC), .D1(VCC), .D2(GND), .E1(VCC),
          .E2(Q), .NS(N_3), .OS(N_2), .OZ(N_1) );
frag_a QL1 ( .A1(J1), .A2(J2NN), .A3(JK), .A4(GND), .A5(J3), .A6(GND), .AZ(N_2) );

endmodule // ttl105q

`endif

`ifdef ttl104q
`else
`define ttl104q
module ttl104q( CLK , CLR, J1, J2, J3, JKNN, K1, K2, K3, PRE, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input PRE /* synthesis syn_isclock=1 */;
input J1, J2, J3, JKNN, K1, K2, K3;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(CLK), .QD(N_2), .QR(CLR), .QS(PRE), .QZ(Q) );
frag_f I_2 ( .F1(K1), .F2(JKNN), .F3(K2), .F4(GND), .F5(K3), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(Q), .B2(GND), .C1(GND), .C2(VCC), .D1(VCC), .D2(GND), .E1(VCC),
          .E2(Q), .NS(N_1), .OS(N_3), .OZ(N_2) );
frag_a QL1 ( .A1(J1), .A2(GND), .A3(J2), .A4(GND), .A5(J3), .A6(JKNN), .AZ(N_3) );

endmodule // ttl104q

`endif

`ifdef ttl08
`else
`define ttl08
module ttl08( A1 , A2, A3, A4, B1, B2, B3, B4, Y1, Y2, Y3, Y4 );
input A1, A2, A3, A4, B1, B2, B3, B4;
output Y1, Y2, Y3, Y4;

and2i0 QL1 ( .A(A4), .B(B4), .Q(Y4) );
and2i0 QL2 ( .A(A3), .B(B3), .Q(Y3) );
and2i0 QL3 ( .A(A2), .B(B2), .Q(Y2) );
and2i0 QL4 ( .A(A1), .B(B1), .Q(Y1) );

endmodule // ttl08

`endif

`ifdef ttl04
`else
`define ttl04
module ttl04( A1 , A2, A3, A4, A5, A6, Y1, Y2, Y3, Y4, Y5, Y6 );
input A1, A2, A3, A4, A5, A6;
output Y1, Y2, Y3, Y4, Y5, Y6;

tri_inv QL1 ( .IN1(A4), .IN2(A5), .IN3(A6), .OUT1(Y4), .OUT2(Y5), .OUT3(Y6) );
tri_inv QL2 ( .IN1(A1), .IN2(A2), .IN3(A3), .OUT1(Y1), .OUT2(Y2), .OUT3(Y3) );

endmodule // ttl04

`endif

`ifdef ttl02
`else
`define ttl02
module ttl02( A1 , A2, A3, A4, B1, B2, B3, B4, Y1, Y2, Y3, Y4 );
input A1, A2, A3, A4, B1, B2, B3, B4;
output Y1, Y2, Y3, Y4;

nor2i0 QL1 ( .A(A2), .B(B2), .Q(Y2) );
nor2i0 QL2 ( .A(A4), .B(B4), .Q(Y4) );
nor2i0 QL3 ( .A(A3), .B(B3), .Q(Y3) );
nor2i0 QL4 ( .A(A1), .B(B1), .Q(Y1) );

endmodule // ttl02

`endif

`ifdef xor5i0
`else
`define xor5i0
module xor5i0( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
supply1 vcc;
supply0 gnd;

logic2 I_5 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(A), .B1(C),
          .B2(gnd), .C1(vcc), .C2(C), .D1(vcc), .D2(C), .E1(C), .E2(gnd),
          .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd), .F5(vcc), .F6(E), .MP(D),
          .MS(E), .NP(D), .NS(E), .OP(B), .OS(A), .OZ(Q), .QC(gnd), .QR(gnd),
          .QS(gnd) );

endmodule // xor5i0

`endif

`ifdef xor4i0
`else
`define xor4i0
module xor4i0( A , B, C, D, Q );
input A, B, C, D;
output Q;
supply1 vcc;
supply0 gnd;

logic2 I_5 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(gnd), .A6(gnd), .B1(C),
          .B2(gnd), .C1(vcc), .C2(C), .D1(vcc), .D2(C), .E1(C), .E2(gnd),
          .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd), .F5(vcc), .F6(B), .MP(D),
          .MS(B), .NP(D), .NS(B), .OP(gnd), .OS(A), .OZ(Q), .QC(gnd), .QR(gnd),
          .QS(gnd) );

endmodule // xor4i0

`endif

`ifdef xor2xor3
`else
`define xor2xor3
module xor2xor3( A0 , A1, B0, B1, C0, Q0, Q1 );
input A0, A1, B0, B1, C0;
output Q0, Q1;
parameter ql_gate = `LOGIC;
supply0 gnd;
supply1 vcc;

lcell2 I_2 ( .A1(gnd), .A2(gnd), .A3(gnd), .A4(gnd), .A5(gnd), .A6(gnd), .B1(B1),
          .B2(gnd), .C1(vcc), .C2(B1), .D1(C0), .D2(gnd), .E1(vcc), .E2(C0),
          .F1(vcc), .F2(B0), .F3(vcc), .F4(gnd), .F5(vcc), .F6(gnd), .MP(gnd),
          .MS(A1), .NP(A0), .NS(B0), .NZ(Q0), .OP(gnd), .OS(gnd), .OZ(Q1),
          .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // xor2xor3

`endif

`ifdef xnor5i0
`else
`define xnor5i0
module xnor5i0( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
supply1 vcc;
supply0 gnd;

logic2 I_5 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(A), .B1(vcc),
          .B2(C), .C1(C), .C2(gnd), .D1(C), .D2(gnd), .E1(vcc), .E2(C), .F1(vcc),
          .F2(gnd), .F3(vcc), .F4(gnd), .F5(vcc), .F6(E), .MP(D), .MS(E), .NP(D),
          .NS(E), .OP(B), .OS(A), .OZ(Q), .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // xnor5i0

`endif

`ifdef xnor4i0
`else
`define xnor4i0
module xnor4i0( A , B, C, D, Q );
input A, B, C, D;
output Q;
supply1 vcc;
supply0 gnd;

logic2 I_5 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(vcc), .B1(vcc),
          .B2(B), .C1(B), .C2(gnd), .D1(B), .D2(gnd), .E1(vcc), .E2(B), .F1(vcc),
          .F2(gnd), .F3(vcc), .F4(gnd), .F5(vcc), .F6(D), .MP(C), .MS(D), .NP(C),
          .NS(D), .OP(gnd), .OS(A), .OZ(Q), .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // xnor4i0

`endif

`ifdef sop16i7
`else
`define sop16i7
module sop16i7( A , B, C, D, E, F, G, H, I, J, K, L, M, N, O, P, Q );
input A, B, C, D, E, F, G, H, I, J, K, L, M, N, O, P;
output Q;
supply1 VCC;
supply0 gnd;

logic2 I_2 ( .A1(A), .A2(D), .A3(B), .A4(E), .A5(C), .A6(F), .B1(H), .B2(I), .C1(VCC),
          .C2(gnd), .D1(VCC), .D2(gnd), .E1(VCC), .E2(gnd), .F1(K), .F2(N),
          .F3(L), .F4(O), .F5(M), .F6(P), .MP(J), .MS(gnd), .NP(J), .NS(gnd),
          .OP(G), .OS(gnd), .OZ(Q), .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // sop16i7

`endif

`ifdef or15i8
`else
`define or15i8
module or15i8( A , B, C, D, E, F, G, H, I, J, K, L, M, N, O, Q );
input A, B, C, D, E, F, G, H, I, J, K, L, M, N, O;
output Q;
supply1 vcc;
supply0 gnd;

logic2 I_2 ( .A1(H), .A2(A), .A3(I), .A4(B), .A5(J), .A6(C), .B1(vcc), .B2(gnd),
          .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd), .E1(D), .E2(gnd), .F1(M),
          .F2(E), .F3(N), .F4(F), .F5(O), .F6(G), .MP(gnd), .MS(gnd), .NP(L),
          .NS(gnd), .OP(K), .OS(gnd), .OZ(Q), .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // or15i8

`endif

`ifdef nor9i5
`else
`define nor9i5
module nor9i5( A , B, C, D, E, F, G, H, I, Q );
input A, B, C, D, E, F, G, H, I;
output Q;
supply0 GND;
supply1 VCC;

logic2 I_1 ( .A1(GND), .A2(GND), .A3(GND), .A4(GND), .A5(GND), .A6(GND), .B1(GND),
          .B2(GND), .C1(GND), .C2(GND), .D1(GND), .D2(GND), .E1(E), .E2(A),
          .F1(G), .F2(B), .F3(H), .F4(C), .F5(I), .F6(D), .MP(GND), .MS(GND),
          .NP(F), .NS(GND), .NZ(Q), .OP(VCC), .OS(GND), .QC(GND), .QR(GND),
          .QS(GND) );

endmodule // nor9i5

`endif

`ifdef nor7i0
`else
`define nor7i0
module nor7i0( A , B, C, D, E, F, G, Q );
input A, B, C, D, E, F, G;
output Q;
supply1 VCC;
supply0 gnd;

logic2 I_2 ( .A1(VCC), .A2(A), .A3(VCC), .A4(B), .A5(VCC), .A6(C), .B1(gnd),
          .B2(gnd), .C1(gnd), .C2(gnd), .D1(gnd), .D2(gnd), .E1(VCC), .E2(D),
          .F1(VCC), .F2(E), .F3(VCC), .F4(F), .F5(VCC), .F6(G), .MP(VCC),
          .MS(gnd), .NP(VCC), .NS(gnd), .OP(VCC), .OS(gnd), .OZ(Q), .QC(gnd),
          .QR(gnd), .QS(gnd) );

endmodule // nor7i0

`endif

`ifdef nor16i9
`else
`define nor16i9
module nor16i9( A , B, C, D, E, F, G, H, I, J, K, L, M, N, O, P, Q );
input A, B, C, D, E, F, G, H, I, J, K, L, M, N, O, P;
output Q;
supply0 gnd;

logic2 I_2 ( .A1(H), .A2(A), .A3(I), .A4(B), .A5(J), .A6(C), .B1(gnd), .B2(gnd),
          .C1(gnd), .C2(gnd), .D1(gnd), .D2(gnd), .E1(L), .E2(D), .F1(N), .F2(E),
          .F3(O), .F4(F), .F5(P), .F6(G), .MP(gnd), .MS(gnd), .NP(M), .NS(gnd),
          .OP(K), .OS(gnd), .OZ(Q), .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // nor16i9

`endif

`ifdef nand8i0
`else
`define nand8i0
module nand8i0( A , B, C, D, E, F, G, H, Q );
input A, B, C, D, E, F, G, H;
output Q;
supply0 GND;
supply1 VCC;

logic2 I_1 ( .A1(A), .A2(GND), .A3(B), .A4(GND), .A5(C), .A6(GND), .B1(VCC),
          .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND), .E2(GND),
          .F1(F), .F2(GND), .F3(G), .F4(GND), .F5(H), .F6(GND), .MP(GND),
          .MS(GND), .NP(E), .NS(GND), .OP(D), .OS(GND), .OZ(Q), .QC(GND),
          .QR(GND), .QS(GND) );

endmodule // nand8i0

`endif

`ifdef nand7i0
`else
`define nand7i0
module nand7i0( A , B, C, D, E, F, G, Q );
input A, B, C, D, E, F, G;
output Q;
supply0 GND;
supply1 VCC;

logic2 I_1 ( .A1(A), .A2(GND), .A3(B), .A4(GND), .A5(C), .A6(GND), .B1(VCC),
          .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND), .E2(GND),
          .F1(F), .F2(GND), .F3(G), .F4(GND), .F5(VCC), .F6(GND), .MP(GND),
          .MS(GND), .NP(E), .NS(GND), .OP(D), .OS(GND), .OZ(Q), .QC(GND),
          .QR(GND), .QS(GND) );

endmodule // nand7i0

`endif

`ifdef nand15i6
`else
`define nand15i6
module nand15i6( A , B, C, D, E, F, G, H, I, J, K, L, M, N, O, Q );
input A, B, C, D, E, F, G, H, I, J, K, L, M, N, O;
output Q;
supply1 vcc;
supply0 gnd;

logic2 I_2 ( .A1(A), .A2(H), .A3(B), .A4(I), .A5(C), .A6(J), .B1(vcc), .B2(gnd),
          .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd), .E1(vcc), .E2(D), .F1(E),
          .F2(M), .F3(F), .F4(N), .F5(G), .F6(O), .MP(gnd), .MS(gnd), .NP(L),
          .NS(gnd), .OP(K), .OS(gnd), .OZ(Q), .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // nand15i6

`endif

`ifdef lshft2q2
`else
`define lshft2q2
module lshft2q2( CLK , CLR, D, Q1, Q2 );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input D;
output Q1, Q2;
wire clk_tst;
wire Qa;
supply1 vcc;
supply0 gnd;

logic2 I_2 ( .A1(gnd), .A2(gnd), .A3(gnd), .A4(gnd), .A5(gnd), .A6(gnd), .B1(Q1),
          .B2(CLR), .C1(Qa), .C2(CLR), .D1(D), .D2(CLR), .E1(Qa), .E2(CLR),
          .F1(CLK), .F2(gnd), .F3(vcc), .F4(gnd), .F5(vcc), .F6(gnd),
          .FZ(clk_tst), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .NZ(Qa),
          .OP(gnd), .OS(gnd), .OZ(Q1), .QC(CLK), .QR(CLR), .QS(gnd), .QZ(Q2) );

endmodule // lshft2q2

`endif

`ifdef logic2
`else
`define logic2
module logic2( A1 , A2, A3, A4, A5, A6, B1, B2, C1, C2, D1, D2, E1, E2, F1, F2,
               F3, F4, F5, F6, MP, MS, NP, NS, OP, OS, QC, QR, QS, AZ, FZ, NZ,
               OZ, QZ );
input A1, A2, A3, A4, A5, A6;
output AZ;
input B1, B2, C1, C2, D1, D2, E1, E2, F1, F2, F3, F4, F5, F6;
output FZ;
input MP, MS, NP, NS;
output NZ;
input OP, OS;
output OZ;
input QC /* synthesis syn_isclock=1 */;
input QR /* synthesis syn_isclock=1 */;
input QS /* synthesis syn_isclock=1 */;
output QZ;
parameter syn_macro = 1, ql_pack = 1;
parameter ql_gate = `LOGIC;

lcell2 I_2 ( .A1(A1), .A2(A2), .A3(A3), .A4(A4), .A5(A5), .A6(A6), .AZ(AZ), .B1(B1),
          .B2(B2), .C1(C1), .C2(C2), .D1(D1), .D2(D2), .E1(E1), .E2(E2), .F1(F1),
          .F2(F2), .F3(F3), .F4(F4), .F5(F5), .F6(F6), .FZ(FZ), .MP(MP), .MS(MS),
          .NP(NP), .NS(NS), .NZ(NZ), .OP(OP), .OS(OS), .OZ(OZ), .QC(QC), .QR(QR),
          .QS(QS), .QZ(QZ) );

endmodule // logic2

`endif

`ifdef ipad8ff
`else
`define ipad8ff
module ipad8ff( FFCLK , FFCLR, FFEN, P, FFQ, Q );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input FFEN;
 output [7:0] FFQ;
 input [7:0] P;
 output [7:0] Q;
parameter syn_macro = 1;

inpadff QL0 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[0]), .P(P[0]),
           .Q(Q[0]) );
inpadff QL1 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[1]), .P(P[1]),
           .Q(Q[1]) );
inpadff QL2 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[2]), .P(P[2]),
           .Q(Q[2]) );
inpadff QL3 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[3]), .P(P[3]),
           .Q(Q[3]) );
inpadff QL4 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[4]), .P(P[4]),
           .Q(Q[4]) );
inpadff QL5 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[5]), .P(P[5]),
           .Q(Q[5]) );
inpadff QL6 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[6]), .P(P[6]),
           .Q(Q[6]) );
inpadff QL7 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[7]), .P(P[7]),
           .Q(Q[7]) );

endmodule // ipad8ff

`endif

`ifdef ipad4ff
`else
`define ipad4ff
module ipad4ff( FFCLK , FFCLR, FFEN, P, FFQ, Q );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input FFEN;
 output [3:0] FFQ;
 input [3:0] P;
 output [3:0] Q;
parameter syn_macro = 1;

inpadff QL0 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[0]), .P(P[0]),
           .Q(Q[0]) );
inpadff QL1 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[1]), .P(P[1]),
           .Q(Q[1]) );
inpadff QL2 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[2]), .P(P[2]),
           .Q(Q[2]) );
inpadff QL3 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[3]), .P(P[3]),
           .Q(Q[3]) );

endmodule // ipad4ff

`endif

`ifdef ipad16ff
`else
`define ipad16ff
module ipad16ff( FFCLK , FFCLR, FFEN, P, FFQ, Q );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input FFEN;
 output [15:0] FFQ;
 input [15:0] P;
 output [15:0] Q;
parameter syn_macro = 1;

inpadff QL0 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[0]), .P(P[0]),
           .Q(Q[0]) );
inpadff QL1 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[1]), .P(P[1]),
           .Q(Q[1]) );
inpadff QL2 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[2]), .P(P[2]),
           .Q(Q[2]) );
inpadff QL3 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[3]), .P(P[3]),
           .Q(Q[3]) );
inpadff QL4 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[4]), .P(P[4]),
           .Q(Q[4]) );
inpadff QL5 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[5]), .P(P[5]),
           .Q(Q[5]) );
inpadff QL6 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[6]), .P(P[6]),
           .Q(Q[6]) );
inpadff QL7 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[7]), .P(P[7]),
           .Q(Q[7]) );
inpadff QL8 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[8]), .P(P[8]),
           .Q(Q[8]) );
inpadff QL9 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[9]), .P(P[9]),
           .Q(Q[9]) );
inpadff QL10 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[10]),
            .P(P[10]), .Q(Q[10]) );
inpadff QL11 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[11]),
            .P(P[11]), .Q(Q[11]) );
inpadff QL12 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[12]),
            .P(P[12]), .Q(Q[12]) );
inpadff QL13 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[13]),
            .P(P[13]), .Q(Q[13]) );
inpadff QL14 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[14]),
            .P(P[14]), .Q(Q[14]) );
inpadff QL15 ( .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN), .FFQ(FFQ[15]),
            .P(P[15]), .Q(Q[15]) );

endmodule // ipad16ff

`endif

`ifdef inpadff
`else
`define inpadff
module inpadff( FFCLK , FFCLR, FFEN, P, FFQ, Q );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input FFEN;
output FFQ;
input P;
output Q;
parameter syn_macro = 1;
parameter ql_gate = `BIDIR;
supply1 VCC;
supply0 GND;

bicell2 QL1 ( .I1(VCC), .I2(GND), .IC(FFCLK), .IE(GND), .IP(P), .IQ(FFQ),
           .IQE(FFEN), .IR(FFCLR), .IZ(Q) );

endmodule // inpadff

`endif

`ifdef hdpadff
`else
`define hdpadff
module hdpadff( FFCLK, FFCLR, FFEN, FFQ, P, Q1 );
input FFCLK /*synthesis syn_isclock=1 */;
input FFCLR /*synthesis syn_isclock=1 */;
input FFEN;
output FFQ;
input P;
output Q1;
parameter syn_macro = 1;
parameter ql_gate = `INCELL;

incell2 QL1 ( .IC(FFCLK), .IP(P), .IQ(FFQ), .IQE(FFEN), .IR(FFCLR), .IZ(Q1) );

endmodule // hdpadff

`endif

`ifdef hdipadff
`else
`define hdipadff
module hdipadff( FFCLK, FFCLR, FFEN, FFQ, P, Q0 );
input FFCLK /*synthesis syn_isclock=1 */;
input FFCLR /*synthesis syn_isclock=1 */;
input FFEN;
output FFQ;
input P;
output Q0;
parameter syn_macro = 1;
parameter ql_gate = `INCELL;

incell2 QL1 ( .IC(FFCLK), .IN(Q0), .IP(P), .IQ(FFQ), .IQE(FFEN), .IR(FFCLR) );

endmodule // hdipadff

`endif

`ifdef hddpadff
`else
`define hddpadff
module hddpadff( FFCLK, FFCLR, FFEN, FFQ, P, Q0, Q1 );
input FFCLK /*synthesis syn_isclock=1 */;
input FFCLR /*synthesis syn_isclock=1 */;
input FFEN;
output FFQ;
input P;
output Q0, Q1;
parameter syn_macro = 1;
parameter ql_gate = `INCELL;

incell2 QL1 ( .IC(FFCLK), .IN(Q0), .IP(P), .IQ(FFQ), .IQE(FFEN), .IR(FFCLR),
           .IZ(Q1) );

endmodule // hddpadff

`endif

`ifdef gclkbuff
`else
`define gclkbuff
module gclkbuff( A , Z );
input A;
output Z;
parameter ql_gate = `HSCK;

bufcell I_1 ( .IC(A), .IZ(Z) );

endmodule // gclkbuff

`endif

`ifdef fstadd8
`else
`define fstadd8
module fstadd8( A , B, CI, SUM );
 input [7:0] A;
 input [7:0] B;
input CI;
 output [7:0] SUM;
wire A3_AND_B3;
wire CI3_N;
wire CI1_N;
wire P1;
wire N_1;
wire P7_N;
wire P5_N;
wire P7;
wire CI7_N;
wire G7;
wire G6;
wire A7_NOR_B7;
wire A6_NOR_B6;
wire P6;
wire CI6_N;
wire CI_6_6;
wire CI_6_4;
wire CI_6_2;
wire G5_N;
wire G5;
wire G4;
wire A5_NOR_B5;
wire A4_NOR_B4;
wire P5;
wire CI5_N;
wire P4;
wire CI4_N;
wire CI_4_4;
wire CI_4_6;
wire CI0_N;
wire CI2_N;
wire P0;
wire P2;
wire CI_2_6;
wire P3;
wire P3_N;
wire P1_N;
wire A0_NOR_B0;
wire A2_NOR_B2;
wire A1_NOR_B1;
wire A3_NOR_B3;
wire G0;
wire G1_N;
wire G1;
wire G2;
wire G3;
supply1 vcc;
supply0 gnd;

logic2 I_54 ( .A1(vcc), .A2(A[2]), .A3(vcc), .A4(gnd), .A5(vcc), .A6(B[2]),
           .B1(vcc), .B2(gnd), .C1(gnd), .C2(gnd), .D1(gnd), .D2(gnd), .E1(gnd),
           .E2(G2), .F1(vcc), .F2(A[3]), .F3(vcc), .F4(B[3]), .F5(vcc), .F6(gnd),
           .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd), .OZ(P3),
           .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_33 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(G1_N), .A6(CI_2_6),
           .AZ(CI3_N), .B1(vcc), .B2(A2_NOR_B2), .C1(A2_NOR_B2), .C2(gnd),
           .D1(G2), .D2(gnd), .E1(vcc), .E2(G2), .F1(vcc), .F2(A3_AND_B3),
           .F3(vcc), .F4(A3_NOR_B3), .F5(vcc), .F6(gnd), .MP(vcc), .MS(gnd),
           .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd), .OZ(SUM[3]), .QC(gnd),
           .QR(gnd), .QS(gnd) );
logic2 I_34 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(CI), .AZ(CI1_N),
           .B1(vcc), .B2(A0_NOR_B0), .C1(A0_NOR_B0), .C2(gnd), .D1(G0),
           .D2(gnd), .E1(vcc), .E2(G0), .F1(vcc), .F2(G1), .F3(vcc),
           .F4(A1_NOR_B1), .F5(vcc), .F6(gnd), .FZ(P1), .MP(vcc), .MS(gnd),
           .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd), .OZ(SUM[1]), .QC(gnd),
           .QR(gnd), .QS(gnd) );
logic2 I_52 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(G1_N), .A5(P3), .A6(gnd),
           .AZ(CI_4_4), .B1(gnd), .B2(gnd), .C1(gnd), .C2(gnd), .D1(gnd),
           .D2(gnd), .E1(P3), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd),
           .F5(CI), .F6(P1_N), .FZ(CI_2_6), .MP(vcc), .MS(gnd), .NP(vcc),
           .NS(gnd), .NZ(CI_4_6), .OP(vcc), .OS(gnd), .QC(gnd), .QR(gnd),
           .QS(gnd) );
logic2 I_53 ( .A1(CI), .A2(P1_N), .A3(P3), .A4(P5_N), .A5(vcc), .A6(gnd),
           .AZ(CI_6_6), .B1(gnd), .B2(gnd), .C1(gnd), .C2(gnd), .D1(gnd),
           .D2(gnd), .E1(vcc), .E2(P5_N), .F1(vcc), .F2(G1_N), .F3(P3),
           .F4(P5_N), .F5(vcc), .F6(gnd), .FZ(CI_6_4), .MP(gnd), .MS(gnd),
           .NP(gnd), .NS(G3), .NZ(CI_6_2), .OP(gnd), .OS(gnd), .QC(gnd),
           .QR(gnd), .QS(gnd) );
logic2 I_48 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(A[6]), .A5(vcc), .A6(B[6]),
           .AZ(A6_NOR_B6), .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc),
           .D2(gnd), .E1(vcc), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(A[7]),
           .F5(vcc), .F6(B[7]), .FZ(A7_NOR_B7), .MP(vcc), .MS(gnd), .NP(vcc),
           .NS(gnd), .OP(vcc), .OS(gnd), .OZ(P7_N), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_51 ( .A1(vcc), .A2(gnd), .A3(A[5]), .A4(gnd), .A5(B[5]), .A6(gnd), .AZ(G5),
           .B1(gnd), .B2(gnd), .C1(B[6]), .C2(gnd), .D1(gnd), .D2(gnd), .E1(gnd),
           .E2(gnd), .F1(A[7]), .F2(gnd), .F3(B[7]), .F4(gnd), .F5(vcc),
           .F6(gnd), .FZ(G7), .MP(gnd), .MS(A[6]), .NP(gnd), .NS(gnd), .OP(gnd),
           .OS(gnd), .OZ(G6), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_49 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(A[4]), .A5(vcc), .A6(B[4]),
           .AZ(A4_NOR_B4), .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc),
           .D2(gnd), .E1(vcc), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(A[5]),
           .F5(vcc), .F6(B[5]), .FZ(A5_NOR_B5), .MP(vcc), .MS(gnd), .NP(vcc),
           .NS(gnd), .OP(vcc), .OS(gnd), .OZ(P5_N), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_50 ( .A1(vcc), .A2(gnd), .A3(A[4]), .A4(gnd), .A5(B[4]), .A6(gnd), .AZ(G4),
           .B1(vcc), .B2(gnd), .C1(vcc), .C2(B[5]), .D1(vcc), .D2(B[5]),
           .E1(gnd), .E2(gnd), .F1(A[5]), .F2(gnd), .F3(B[5]), .F4(gnd),
           .F5(vcc), .F6(gnd), .FZ(N_1), .MP(gnd), .MS(A[5]), .NP(gnd),
           .NS(A[5]), .OP(vcc), .OS(gnd), .OZ(G5_N), .QC(gnd), .QR(gnd),
           .QS(gnd) );
logic2 I_44 ( .A1(vcc), .A2(G3), .A3(vcc), .A4(CI_4_4), .A5(vcc), .A6(CI_4_6),
           .AZ(CI5_N), .B1(vcc), .B2(A4_NOR_B4), .C1(A4_NOR_B4), .C2(gnd),
           .D1(G4), .D2(gnd), .E1(vcc), .E2(G4), .F1(vcc), .F2(G5), .F3(vcc),
           .F4(A5_NOR_B5), .F5(vcc), .F6(gnd), .FZ(P5), .MP(vcc), .MS(gnd),
           .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd), .OZ(SUM[5]), .QC(gnd),
           .QR(gnd), .QS(gnd) );
logic2 I_45 ( .A1(G5_N), .A2(CI_6_2), .A3(vcc), .A4(CI_6_4), .A5(vcc), .A6(CI_6_6),
           .AZ(CI7_N), .B1(vcc), .B2(A6_NOR_B6), .C1(A6_NOR_B6), .C2(gnd),
           .D1(G6), .D2(gnd), .E1(vcc), .E2(G6), .F1(vcc), .F2(G7), .F3(vcc),
           .F4(A7_NOR_B7), .F5(vcc), .F6(gnd), .FZ(P7), .MP(vcc), .MS(gnd),
           .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd), .OZ(SUM[7]), .QC(gnd),
           .QR(gnd), .QS(gnd) );
logic2 I_46 ( .A1(vcc), .A2(G3), .A3(vcc), .A4(CI_4_4), .A5(vcc), .A6(CI_4_6),
           .AZ(CI4_N), .B1(vcc), .B2(B[4]), .C1(B[4]), .C2(gnd), .D1(B[4]),
           .D2(gnd), .E1(vcc), .E2(B[4]), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd),
           .F5(gnd), .F6(gnd), .MP(gnd), .MS(A[4]), .NP(gnd), .NS(A[4]), .NZ(P4),
           .OP(vcc), .OS(gnd), .OZ(SUM[4]), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_47 ( .A1(G5_N), .A2(CI_6_2), .A3(vcc), .A4(CI_6_4), .A5(vcc), .A6(CI_6_6),
           .AZ(CI6_N), .B1(vcc), .B2(B[6]), .C1(B[6]), .C2(gnd), .D1(B[6]),
           .D2(gnd), .E1(vcc), .E2(B[6]), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd),
           .F5(vcc), .F6(gnd), .MP(gnd), .MS(A[6]), .NP(gnd), .NS(A[6]), .NZ(P6),
           .OP(vcc), .OS(gnd), .OZ(SUM[6]), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_23 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(CI), .AZ(CI0_N),
           .B1(vcc), .B2(B[0]), .C1(B[0]), .C2(gnd), .D1(B[0]), .D2(gnd),
           .E1(vcc), .E2(B[0]), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd), .F5(gnd),
           .F6(gnd), .MP(gnd), .MS(A[0]), .NP(gnd), .NS(A[0]), .NZ(P0), .OP(vcc),
           .OS(gnd), .OZ(SUM[0]), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_21 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(G1_N), .A6(CI_2_6),
           .AZ(CI2_N), .B1(vcc), .B2(B[2]), .C1(B[2]), .C2(gnd), .D1(B[2]),
           .D2(gnd), .E1(vcc), .E2(B[2]), .F1(A[3]), .F2(gnd), .F3(B[3]),
           .F4(gnd), .F5(vcc), .F6(gnd), .FZ(A3_AND_B3), .MP(gnd), .MS(A[2]),
           .NP(gnd), .NS(A[2]), .NZ(P2), .OP(vcc), .OS(gnd), .OZ(SUM[2]),
           .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_37 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(A[2]), .A5(vcc), .A6(B[2]),
           .AZ(A2_NOR_B2), .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc),
           .D2(gnd), .E1(vcc), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(A[3]),
           .F5(vcc), .F6(B[3]), .FZ(A3_NOR_B3), .MP(vcc), .MS(gnd), .NP(vcc),
           .NS(gnd), .OP(vcc), .OS(gnd), .OZ(P3_N), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_36 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(A[0]), .A5(vcc), .A6(B[0]),
           .AZ(A0_NOR_B0), .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc),
           .D2(gnd), .E1(vcc), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(A[1]),
           .F5(vcc), .F6(B[1]), .FZ(A1_NOR_B1), .MP(vcc), .MS(gnd), .NP(vcc),
           .NS(gnd), .OP(vcc), .OS(gnd), .OZ(P1_N), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_6 ( .A1(vcc), .A2(gnd), .A3(A[0]), .A4(gnd), .A5(B[0]), .A6(gnd), .AZ(G0),
          .B1(vcc), .B2(gnd), .C1(vcc), .C2(B[1]), .D1(vcc), .D2(B[1]), .E1(gnd),
          .E2(gnd), .F1(A[1]), .F2(gnd), .F3(B[1]), .F4(gnd), .F5(vcc), .F6(gnd),
          .FZ(G1), .MP(gnd), .MS(A[1]), .NP(gnd), .NS(A[1]), .OP(vcc), .OS(gnd),
          .OZ(G1_N), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_12 ( .A1(vcc), .A2(gnd), .A3(A[2]), .A4(gnd), .A5(B[2]), .A6(gnd), .AZ(G2),
           .B1(gnd), .B2(gnd), .C1(B[3]), .C2(gnd), .D1(B[3]), .D2(gnd),
           .E1(vcc), .E2(gnd), .F1(A[3]), .F2(gnd), .F3(B[3]), .F4(gnd),
           .F5(vcc), .F6(gnd), .MP(gnd), .MS(A[3]), .NP(gnd), .NS(A[3]),
           .OP(vcc), .OS(gnd), .OZ(G3), .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // fstadd8

`endif

`ifdef fstadd4
`else
`define fstadd4
module fstadd4( A , B, CI, SUM );
 input [3:0] A;
 input [3:0] B;
input CI;
 output [3:0] SUM;
wire CI_2_6;
wire P1_N;
wire CI0_N;
wire CI2_N;
wire CI1_N;
wire CI3_N;
wire A0_NOR_B0;
wire A2_NOR_B2;
wire A1_NOR_B1;
wire A3_NOR_B3;
wire G0;
wire G1_N;
wire G1;
wire G2;
wire G3;
supply1 vcc;
supply0 gnd;

logic2 I_23 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(CI), .AZ(CI0_N),
           .B1(vcc), .B2(B[0]), .C1(B[0]), .C2(gnd), .D1(B[0]), .D2(gnd),
           .E1(vcc), .E2(B[0]), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd), .F5(gnd),
           .F6(gnd), .MP(gnd), .MS(A[0]), .NP(gnd), .NS(A[0]), .OP(vcc),
           .OS(gnd), .OZ(SUM[0]), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_21 ( .A1(vcc), .A2(gnd), .A3(G1_N), .A4(gnd), .A5(vcc), .A6(CI_2_6),
           .AZ(CI2_N), .B1(vcc), .B2(B[2]), .C1(B[2]), .C2(gnd), .D1(B[2]),
           .D2(gnd), .E1(vcc), .E2(B[2]), .F1(CI), .F2(P1_N), .F3(vcc), .F4(gnd),
           .F5(vcc), .F6(gnd), .FZ(CI_2_6), .MP(gnd), .MS(A[2]), .NP(gnd),
           .NS(A[2]), .OP(vcc), .OS(gnd), .OZ(SUM[2]), .QC(gnd), .QR(gnd),
           .QS(gnd) );
logic2 I_37 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(A[2]), .A5(vcc), .A6(B[2]),
           .AZ(A2_NOR_B2), .B1(gnd), .B2(gnd), .C1(B[2]), .C2(gnd), .D1(gnd),
           .D2(gnd), .E1(A[3]), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc),
           .F4(A[3]), .F5(vcc), .F6(B[3]), .FZ(A3_NOR_B3), .MP(gnd), .MS(A[2]),
           .NP(gnd), .NS(B[3]), .NZ(G3), .OP(gnd), .OS(gnd), .OZ(G2), .QC(gnd),
           .QR(gnd), .QS(gnd) );
logic2 I_33 ( .A1(vcc), .A2(gnd), .A3(G1_N), .A4(gnd), .A5(vcc), .A6(CI_2_6),
           .AZ(CI3_N), .B1(vcc), .B2(A2_NOR_B2), .C1(A2_NOR_B2), .C2(gnd),
           .D1(G2), .D2(gnd), .E1(vcc), .E2(G2), .F1(vcc), .F2(G3), .F3(vcc),
           .F4(A3_NOR_B3), .F5(vcc), .F6(gnd), .MP(vcc), .MS(gnd), .NP(vcc),
           .NS(gnd), .OP(vcc), .OS(gnd), .OZ(SUM[3]), .QC(gnd), .QR(gnd),
           .QS(gnd) );
logic2 I_34 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(CI), .AZ(CI1_N),
           .B1(vcc), .B2(A0_NOR_B0), .C1(A0_NOR_B0), .C2(gnd), .D1(G0),
           .D2(gnd), .E1(vcc), .E2(G0), .F1(vcc), .F2(G1), .F3(vcc),
           .F4(A1_NOR_B1), .F5(vcc), .F6(gnd), .MP(vcc), .MS(gnd), .NP(vcc),
           .NS(gnd), .OP(vcc), .OS(gnd), .OZ(SUM[1]), .QC(gnd), .QR(gnd),
           .QS(gnd) );
logic2 I_6 ( .A1(vcc), .A2(gnd), .A3(A[0]), .A4(gnd), .A5(B[0]), .A6(gnd), .AZ(G0),
          .B1(vcc), .B2(gnd), .C1(vcc), .C2(B[1]), .D1(vcc), .D2(B[1]), .E1(gnd),
          .E2(gnd), .F1(A[1]), .F2(gnd), .F3(B[1]), .F4(gnd), .F5(vcc), .F6(gnd),
          .FZ(G1), .MP(gnd), .MS(A[1]), .NP(gnd), .NS(A[1]), .OP(vcc), .OS(gnd),
          .OZ(G1_N), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_12 ( .A1(vcc), .A2(A[0]), .A3(vcc), .A4(B[0]), .A5(vcc), .A6(gnd),
           .AZ(A0_NOR_B0), .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc),
           .D2(gnd), .E1(vcc), .E2(gnd), .F1(vcc), .F2(A[1]), .F3(vcc),
           .F4(B[1]), .F5(vcc), .F6(gnd), .FZ(A1_NOR_B1), .MP(vcc), .MS(gnd),
           .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd), .OZ(P1_N), .QC(gnd), .QR(gnd),
           .QS(gnd) );

endmodule // fstadd4

`endif

`ifdef fstadd16
`else
`define fstadd16
module fstadd16( A , B, CI, SUM );
 input [15:0] A;
 input [15:0] B;
input CI;
 output [15:0] SUM;
wire G15;
wire A7_AND_B7;
wire N_4;
wire A7_XOR_B7;
wire CI14_N;
wire A15_AND_B15;
wire A9_XOR_B9;
wire P15_N;
wire P13_N;
wire T1_12_6;
wire P15;
wire P13;
wire G11;
wire P11;
wire P11_N;
wire CI_16_3;
wire CI_16_5;
wire CI_16_6;
wire CI15_N;
wire G14;
wire A15_NOR_B15;
wire A14_NOR_B14;
wire A15_XOR_B15;
wire G13_N;
wire CI_14_2;
wire CI_14_3;
wire CI_14_4;
wire CI_14_5;
wire CI_14_6;
wire CI10_N;
wire P10;
wire CI11_N;
wire A10_NOR_B10;
wire A10_AND_B10;
wire A11_XOR_B11;
wire A11_NOR_B11;
wire CI12_N;
wire P12;
wire CI_12_1;
wire CI_12_2;
wire CI_12_3;
wire CI_12_4;
wire CI_12_6;
wire CI13_N;
wire A12_NOR_B12;
wire G12;
wire A13_XOR_B13;
wire G13;
wire A13_NOR_B13;
wire CI4_N;
wire CI6_N;
wire P4;
wire P6;
wire A11_AND_B11;
wire CI5_N;
wire CI7_N;
wire P5;
wire G9_N;
wire P7_N;
wire CI_10_3;
wire CI_10_5;
wire CI_10_6;
wire CI_10_2;
wire P9_N;
wire CI_10_4;
wire P9;
wire CI9_N;
wire A9_NOR_B9;
wire G9;
wire G8;
wire A8_NOR_B8;
wire CI8_N;
wire P8;
wire CI_8_6;
wire CI_8_5;
wire CI_8_4;
wire CI_8_3;
wire P7;
wire A3_AND_B3;
wire CI3_N;
wire CI1_N;
wire P1;
wire P5_N;
wire G7;
wire G6;
wire A7_NOR_B7;
wire A6_NOR_B6;
wire CI_6_6;
wire CI_6_4;
wire CI_6_2;
wire G5_N;
wire G5;
wire G4;
wire A5_NOR_B5;
wire A4_NOR_B4;
wire CI_4_4;
wire CI_4_6;
wire CI0_N;
wire CI2_N;
wire P0;
wire P2;
wire CI_2_6;
wire P3;
wire P3_N;
wire P1_N;
wire A0_NOR_B0;
wire A2_NOR_B2;
wire A1_NOR_B1;
wire A3_NOR_B3;
wire G0;
wire G1_N;
wire G1;
wire G2;
wire G3;
supply1 vcc;
supply0 gnd;

logic2 I_106 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(A[6]), .A5(vcc), .A6(B[6]),
            .B1(vcc), .B2(gnd), .C1(gnd), .C2(gnd), .D1(gnd), .D2(gnd), .E1(gnd),
            .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(A[7]), .F5(vcc),
            .F6(B[7]), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc),
            .OS(gnd), .OZ(P7), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_99 ( .A1(vcc), .A2(gnd), .A3(A[14]), .A4(gnd), .A5(B[14]), .A6(gnd),
           .AZ(G14), .B1(vcc), .B2(gnd), .C1(B[15]), .C2(gnd), .D1(B[15]),
           .D2(gnd), .E1(vcc), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd),
           .F5(vcc), .F6(gnd), .MP(gnd), .MS(A[15]), .NP(gnd), .NS(A[15]),
           .OP(vcc), .OS(gnd), .OZ(G15), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_81 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(A[10]), .A5(vcc), .A6(B[10]),
           .AZ(N_4), .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd),
           .E1(vcc), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(A[11]),
           .F5(vcc), .F6(B[11]), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd),
           .OP(vcc), .OS(gnd), .OZ(P11_N), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_96 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(P7), .A6(G5_N), .B1(gnd),
           .B2(gnd), .C1(G7), .C2(gnd), .D1(gnd), .D2(gnd), .E1(vcc), .E2(gnd),
           .F1(vcc), .F2(P11_N), .F3(P9), .F4(P13_N), .F5(vcc), .F6(gnd),
           .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd),
           .OZ(CI_14_4), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_84 ( .A1(vcc), .A2(gnd), .A3(A[10]), .A4(gnd), .A5(B[10]), .A6(gnd),
           .AZ(A10_AND_B10), .B1(gnd), .B2(gnd), .C1(B[11]), .C2(gnd),
           .D1(B[11]), .D2(gnd), .E1(vcc), .E2(gnd), .F1(vcc), .F2(gnd),
           .F3(A[13]), .F4(gnd), .F5(B[13]), .F6(gnd), .FZ(G13), .MP(gnd),
           .MS(A[11]), .NP(gnd), .NS(A[11]), .OP(vcc), .OS(gnd), .OZ(G11),
           .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_97 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(B[14]), .A5(vcc), .A6(A[14]),
           .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd), .E1(vcc),
           .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(B[15]), .F5(vcc),
           .F6(A[15]), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc),
           .OS(gnd), .OZ(P15_N), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_98 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(B[14]), .A5(vcc), .A6(A[14]),
           .AZ(A14_NOR_B14), .B1(vcc), .B2(gnd), .C1(gnd), .C2(gnd), .D1(gnd),
           .D2(gnd), .E1(gnd), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc),
           .F4(B[15]), .F5(vcc), .F6(A[15]), .FZ(A15_NOR_B15), .MP(vcc),
           .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd), .OZ(P15), .QC(gnd),
           .QR(gnd), .QS(gnd) );
logic2 I_92 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(A[12]), .A5(vcc), .A6(B[12]),
           .AZ(A12_NOR_B12), .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc),
           .D2(gnd), .E1(vcc), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc),
           .F4(A[13]), .F5(vcc), .F6(B[13]), .FZ(A13_NOR_B13), .MP(vcc),
           .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd), .OZ(P13_N),
           .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_93 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(A[12]), .A5(vcc), .A6(B[12]),
           .B1(vcc), .B2(gnd), .C1(gnd), .C2(gnd), .D1(gnd), .D2(gnd), .E1(gnd),
           .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(A[13]), .F5(vcc),
           .F6(B[13]), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc),
           .OS(gnd), .OZ(P13), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_95 ( .A1(vcc), .A2(G9_N), .A3(vcc), .A4(P11_N), .A5(vcc), .A6(gnd),
           .B1(gnd), .B2(gnd), .C1(G11), .C2(gnd), .D1(gnd), .D2(gnd), .E1(vcc),
           .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd), .F5(vcc),
           .F6(P13_N), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc),
           .OS(gnd), .OZ(CI_14_2), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_85 ( .A1(G11), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(gnd), .B1(vcc),
           .B2(gnd), .C1(gnd), .C2(gnd), .D1(gnd), .D2(gnd), .E1(gnd), .E2(gnd),
           .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd), .F5(P11), .F6(G9_N), .MP(vcc),
           .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd), .OZ(CI_12_1),
           .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_86 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(P15), .A6(gnd), .B1(vcc),
           .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd), .E1(vcc), .E2(P13),
           .F1(vcc), .F2(P5_N), .F3(G3), .F4(P7_N), .F5(P9), .F6(P11_N),
           .FZ(CI_12_2), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .NZ(CI_14_3),
           .OP(vcc), .OS(gnd), .OZ(CI_16_3), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_82 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(A[10]), .A5(vcc), .A6(B[10]),
           .AZ(A10_NOR_B10), .B1(vcc), .B2(gnd), .C1(gnd), .C2(gnd), .D1(gnd),
           .D2(gnd), .E1(gnd), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc),
           .F4(A[11]), .F5(vcc), .F6(B[11]), .FZ(A11_NOR_B11), .MP(vcc),
           .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd), .OZ(P11), .QC(gnd),
           .QR(gnd), .QS(gnd) );
logic2 I_90 ( .A1(P15), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(gnd), .B1(gnd),
           .B2(gnd), .C1(gnd), .C2(gnd), .D1(gnd), .D2(gnd), .E1(P13), .E2(gnd),
           .F1(P11), .F2(P7_N), .F3(P9), .F4(P5_N), .F5(P3), .F6(T1_12_6),
           .FZ(CI_12_6), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .NZ(CI_14_6),
           .OP(vcc), .OS(gnd), .OZ(CI_16_6), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_91 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(B[0]), .A5(vcc), .A6(A[0]),
           .B1(vcc), .B2(CI), .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd), .E1(vcc),
           .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(B[1]), .F5(vcc),
           .F6(A[1]), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd),
           .OZ(T1_12_6), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_88 ( .A1(vcc), .A2(G5_N), .A3(vcc), .A4(P7_N), .A5(vcc), .A6(gnd),
           .B1(vcc), .B2(gnd), .C1(vcc), .C2(G7), .D1(vcc), .D2(gnd), .E1(gnd),
           .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd), .F5(P9), .F6(P11_N),
           .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd),
           .OZ(CI_12_3), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_89 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(P15), .A6(gnd), .B1(vcc),
           .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd), .E1(vcc), .E2(P13),
           .F1(P11), .F2(P7_N), .F3(P9), .F4(P5_N), .F5(P3), .F6(G1_N),
           .FZ(CI_12_4), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .NZ(CI_14_5),
           .OP(vcc), .OS(gnd), .OZ(CI_16_5), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_66 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(A[8]), .A5(vcc), .A6(B[8]),
           .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd), .E1(vcc),
           .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(A[9]), .F5(vcc),
           .F6(B[9]), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd),
           .OZ(P9_N), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_67 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(A[8]), .A5(vcc), .A6(B[8]),
           .B1(vcc), .B2(gnd), .C1(gnd), .C2(gnd), .D1(gnd), .D2(gnd), .E1(gnd),
           .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(A[9]), .F5(vcc),
           .F6(B[9]), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd),
           .OZ(P9), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_83 ( .A1(vcc), .A2(gnd), .A3(A[12]), .A4(gnd), .A5(B[12]), .A6(gnd),
           .AZ(G12), .B1(vcc), .B2(gnd), .C1(vcc), .C2(B[13]), .D1(vcc),
           .D2(B[13]), .E1(gnd), .E2(gnd), .F1(vcc), .F2(gnd), .F3(A[15]),
           .F4(gnd), .F5(B[15]), .F6(gnd), .FZ(A15_AND_B15), .MP(gnd),
           .MS(A[13]), .NP(gnd), .NS(A[13]), .OP(vcc), .OS(gnd), .OZ(G13_N),
           .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_50 ( .A1(vcc), .A2(gnd), .A3(A[4]), .A4(gnd), .A5(B[4]), .A6(gnd), .AZ(G4),
           .B1(vcc), .B2(gnd), .C1(vcc), .C2(B[5]), .D1(vcc), .D2(B[5]),
           .E1(gnd), .E2(gnd), .F1(A[7]), .F2(gnd), .F3(B[7]), .F4(gnd),
           .F5(vcc), .F6(gnd), .FZ(A7_AND_B7), .MP(gnd), .MS(A[5]), .NP(gnd),
           .NS(A[5]), .OP(vcc), .OS(gnd), .OZ(G5_N), .QC(gnd), .QR(gnd),
           .QS(gnd) );
logic2 I_76 ( .A1(G13_N), .A2(CI_14_2), .A3(CI_14_3), .A4(CI_14_4), .A5(CI_14_5),
           .A6(CI_14_6), .AZ(CI15_N), .B1(vcc), .B2(A14_NOR_B14),
           .C1(A14_NOR_B14), .C2(gnd), .D1(G14), .D2(gnd), .E1(vcc), .E2(G14),
           .F1(vcc), .F2(A15_AND_B15), .F3(vcc), .F4(A15_NOR_B15), .F5(vcc),
           .F6(gnd), .FZ(A15_XOR_B15), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd),
           .OP(vcc), .OS(gnd), .OZ(SUM[15]), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_77 ( .A1(G13_N), .A2(CI_14_2), .A3(CI_14_3), .A4(CI_14_4), .A5(CI_14_5),
           .A6(CI_14_6), .AZ(CI14_N), .B1(vcc), .B2(A[14]), .C1(A[14]),
           .C2(gnd), .D1(A[14]), .D2(gnd), .E1(vcc), .E2(A[14]), .F1(vcc),
           .F2(gnd), .F3(vcc), .F4(gnd), .F5(gnd), .F6(gnd), .MP(gnd),
           .MS(B[14]), .NP(gnd), .NS(B[14]), .OP(vcc), .OS(gnd), .OZ(SUM[14]),
           .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_71 ( .A1(G9_N), .A2(CI_10_2), .A3(CI_10_3), .A4(CI_10_4), .A5(CI_10_5),
           .A6(CI_10_6), .AZ(CI11_N), .B1(vcc), .B2(A10_NOR_B10),
           .C1(A10_NOR_B10), .C2(gnd), .D1(A10_AND_B10), .D2(gnd), .E1(vcc),
           .E2(A10_AND_B10), .F1(vcc), .F2(A11_AND_B11), .F3(vcc),
           .F4(A11_NOR_B11), .F5(vcc), .F6(gnd), .FZ(A11_XOR_B11), .MP(vcc),
           .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd), .OZ(SUM[11]),
           .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_72 ( .A1(G9_N), .A2(CI_10_2), .A3(CI_10_3), .A4(CI_10_4), .A5(CI_10_5),
           .A6(CI_10_6), .AZ(CI10_N), .B1(vcc), .B2(A[10]), .C1(A[10]),
           .C2(gnd), .D1(A[10]), .D2(gnd), .E1(vcc), .E2(A[10]), .F1(vcc),
           .F2(gnd), .F3(vcc), .F4(A[9]), .F5(vcc), .F6(B[9]), .FZ(A9_NOR_B9),
           .MP(gnd), .MS(B[10]), .NP(gnd), .NS(B[10]), .NZ(P10), .OP(vcc),
           .OS(gnd), .OZ(SUM[10]), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_75 ( .A1(CI_12_1), .A2(CI_12_2), .A3(CI_12_3), .A4(CI_12_4), .A5(vcc),
           .A6(CI_12_6), .AZ(CI12_N), .B1(vcc), .B2(A[12]), .C1(A[12]),
           .C2(gnd), .D1(A[12]), .D2(gnd), .E1(vcc), .E2(A[12]), .F1(vcc),
           .F2(gnd), .F3(vcc), .F4(A[8]), .F5(vcc), .F6(B[8]), .FZ(A8_NOR_B8),
           .MP(gnd), .MS(B[12]), .NP(gnd), .NS(B[12]), .NZ(P12), .OP(vcc),
           .OS(gnd), .OZ(SUM[12]), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_74 ( .A1(CI_12_1), .A2(CI_12_2), .A3(CI_12_3), .A4(CI_12_4), .A5(vcc),
           .A6(CI_12_6), .AZ(CI13_N), .B1(vcc), .B2(A12_NOR_B12),
           .C1(A12_NOR_B12), .C2(gnd), .D1(G12), .D2(gnd), .E1(vcc), .E2(G12),
           .F1(vcc), .F2(G13), .F3(vcc), .F4(A13_NOR_B13), .F5(vcc), .F6(gnd),
           .FZ(A13_XOR_B13), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc),
           .OS(gnd), .OZ(SUM[13]), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_45 ( .A1(G5_N), .A2(CI_6_2), .A3(vcc), .A4(CI_6_4), .A5(vcc), .A6(CI_6_6),
           .AZ(CI7_N), .B1(vcc), .B2(A6_NOR_B6), .C1(A6_NOR_B6), .C2(gnd),
           .D1(G6), .D2(gnd), .E1(vcc), .E2(G6), .F1(vcc), .F2(A7_AND_B7),
           .F3(vcc), .F4(A7_NOR_B7), .F5(vcc), .F6(gnd), .FZ(A7_XOR_B7),
           .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd),
           .OZ(SUM[7]), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_47 ( .A1(G5_N), .A2(CI_6_2), .A3(vcc), .A4(CI_6_4), .A5(vcc), .A6(CI_6_6),
           .AZ(CI6_N), .B1(vcc), .B2(B[6]), .C1(B[6]), .C2(gnd), .D1(B[6]),
           .D2(gnd), .E1(vcc), .E2(B[6]), .F1(vcc), .F2(gnd), .F3(A[11]),
           .F4(gnd), .F5(B[11]), .F6(gnd), .FZ(A11_AND_B11), .MP(gnd),
           .MS(A[6]), .NP(gnd), .NS(A[6]), .NZ(P6), .OP(vcc), .OS(gnd),
           .OZ(SUM[6]), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_44 ( .A1(vcc), .A2(G3), .A3(vcc), .A4(CI_4_4), .A5(vcc), .A6(CI_4_6),
           .AZ(CI5_N), .B1(vcc), .B2(A4_NOR_B4), .C1(A4_NOR_B4), .C2(gnd),
           .D1(G4), .D2(gnd), .E1(vcc), .E2(G4), .F1(vcc), .F2(G5), .F3(vcc),
           .F4(A5_NOR_B5), .F5(vcc), .F6(gnd), .FZ(P5), .MP(vcc), .MS(gnd),
           .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd), .OZ(SUM[5]), .QC(gnd),
           .QR(gnd), .QS(gnd) );
logic2 I_46 ( .A1(vcc), .A2(G3), .A3(vcc), .A4(CI_4_4), .A5(vcc), .A6(CI_4_6),
           .AZ(CI4_N), .B1(vcc), .B2(B[4]), .C1(B[4]), .C2(gnd), .D1(B[4]),
           .D2(gnd), .E1(vcc), .E2(B[4]), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd),
           .F5(gnd), .F6(gnd), .MP(gnd), .MS(A[4]), .NP(gnd), .NS(A[4]), .NZ(P4),
           .OP(vcc), .OS(gnd), .OZ(SUM[4]), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_68 ( .A1(vcc), .A2(gnd), .A3(A[8]), .A4(gnd), .A5(B[8]), .A6(gnd), .AZ(G8),
           .B1(vcc), .B2(gnd), .C1(vcc), .C2(B[9]), .D1(vcc), .D2(B[9]),
           .E1(gnd), .E2(gnd), .F1(A[9]), .F2(gnd), .F3(B[9]), .F4(gnd),
           .F5(vcc), .F6(gnd), .FZ(G9), .MP(gnd), .MS(A[9]), .NP(gnd), .NS(A[9]),
           .OP(vcc), .OS(gnd), .OZ(G9_N), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_6 ( .A1(vcc), .A2(gnd), .A3(A[0]), .A4(gnd), .A5(B[0]), .A6(gnd), .AZ(G0),
          .B1(vcc), .B2(gnd), .C1(vcc), .C2(B[1]), .D1(vcc), .D2(B[1]), .E1(gnd),
          .E2(gnd), .F1(A[1]), .F2(gnd), .F3(B[1]), .F4(gnd), .F5(vcc), .F6(gnd),
          .FZ(G1), .MP(gnd), .MS(A[1]), .NP(gnd), .NS(A[1]), .OP(vcc), .OS(gnd),
          .OZ(G1_N), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_48 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(A[6]), .A5(vcc), .A6(B[6]),
           .AZ(A6_NOR_B6), .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc),
           .D2(gnd), .E1(vcc), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(A[7]),
           .F5(vcc), .F6(B[7]), .FZ(A7_NOR_B7), .MP(vcc), .MS(gnd), .NP(vcc),
           .NS(gnd), .OP(vcc), .OS(gnd), .OZ(P7_N), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_65 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(P9_N), .B1(vcc),
           .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd), .E1(vcc), .E2(P7),
           .F1(vcc), .F2(gnd), .F3(vcc), .F4(G1_N), .F5(P3), .F6(P5_N),
           .FZ(CI_6_4), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .NZ(CI_8_5),
           .OP(vcc), .OS(gnd), .OZ(CI_10_5), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_64 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(P9_N), .B1(vcc),
           .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd), .E1(vcc), .E2(P7),
           .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd), .F5(G3), .F6(P5_N),
           .FZ(CI_6_2), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .NZ(CI_8_3),
           .OP(vcc), .OS(gnd), .OZ(CI_10_3), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_62 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(P9_N), .B1(gnd),
           .B2(gnd), .C1(gnd), .C2(gnd), .D1(gnd), .D2(gnd), .E1(P7), .E2(gnd),
           .F1(vcc), .F2(gnd), .F3(CI), .F4(P1_N), .F5(P3), .F6(P5_N),
           .FZ(CI_6_6), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .NZ(CI_8_6),
           .OP(vcc), .OS(gnd), .OZ(CI_10_6), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_60 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(G7), .A6(P9_N),
           .AZ(CI_10_2), .B1(gnd), .B2(gnd), .C1(gnd), .C2(gnd), .D1(gnd),
           .D2(gnd), .E1(vcc), .E2(P9_N), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd),
           .F5(P7), .F6(G5_N), .FZ(CI_8_4), .MP(vcc), .MS(gnd), .NP(vcc),
           .NS(gnd), .NZ(CI_10_4), .OP(vcc), .OS(gnd), .QC(gnd), .QR(gnd),
           .QS(gnd) );
logic2 I_58 ( .A1(vcc), .A2(G7), .A3(CI_8_3), .A4(CI_8_4), .A5(CI_8_5),
           .A6(CI_8_6), .AZ(CI9_N), .B1(vcc), .B2(A8_NOR_B8), .C1(A8_NOR_B8),
           .C2(gnd), .D1(G8), .D2(gnd), .E1(vcc), .E2(G8), .F1(vcc), .F2(G9),
           .F3(vcc), .F4(A9_NOR_B9), .F5(vcc), .F6(gnd), .FZ(A9_XOR_B9),
           .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd),
           .OZ(SUM[9]), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_59 ( .A1(vcc), .A2(G7), .A3(CI_8_3), .A4(CI_8_4), .A5(CI_8_5),
           .A6(CI_8_6), .AZ(CI8_N), .B1(vcc), .B2(B[8]), .C1(B[8]), .C2(gnd),
           .D1(B[8]), .D2(gnd), .E1(vcc), .E2(B[8]), .F1(vcc), .F2(gnd),
           .F3(vcc), .F4(gnd), .F5(vcc), .F6(gnd), .MP(gnd), .MS(A[8]), .NP(gnd),
           .NS(A[8]), .NZ(P8), .OP(vcc), .OS(gnd), .OZ(SUM[8]), .QC(gnd),
           .QR(gnd), .QS(gnd) );
logic2 I_54 ( .A1(vcc), .A2(A[2]), .A3(vcc), .A4(gnd), .A5(vcc), .A6(B[2]),
           .B1(vcc), .B2(gnd), .C1(gnd), .C2(gnd), .D1(gnd), .D2(gnd), .E1(gnd),
           .E2(gnd), .F1(vcc), .F2(A[3]), .F3(vcc), .F4(B[3]), .F5(vcc),
           .F6(gnd), .MP(vcc), .MS(gnd), .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd),
           .OZ(P3), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_33 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(G1_N), .A6(CI_2_6),
           .AZ(CI3_N), .B1(vcc), .B2(A2_NOR_B2), .C1(A2_NOR_B2), .C2(gnd),
           .D1(G2), .D2(gnd), .E1(vcc), .E2(G2), .F1(vcc), .F2(A3_AND_B3),
           .F3(vcc), .F4(A3_NOR_B3), .F5(vcc), .F6(gnd), .MP(vcc), .MS(gnd),
           .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd), .OZ(SUM[3]), .QC(gnd),
           .QR(gnd), .QS(gnd) );
logic2 I_34 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(CI), .AZ(CI1_N),
           .B1(vcc), .B2(A0_NOR_B0), .C1(A0_NOR_B0), .C2(gnd), .D1(G0),
           .D2(gnd), .E1(vcc), .E2(G0), .F1(vcc), .F2(G1), .F3(vcc),
           .F4(A1_NOR_B1), .F5(vcc), .F6(gnd), .FZ(P1), .MP(vcc), .MS(gnd),
           .NP(vcc), .NS(gnd), .OP(vcc), .OS(gnd), .OZ(SUM[1]), .QC(gnd),
           .QR(gnd), .QS(gnd) );
logic2 I_52 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(G1_N), .A5(P3), .A6(gnd),
           .AZ(CI_4_4), .B1(gnd), .B2(gnd), .C1(gnd), .C2(gnd), .D1(gnd),
           .D2(gnd), .E1(P3), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd),
           .F5(CI), .F6(P1_N), .FZ(CI_2_6), .MP(vcc), .MS(gnd), .NP(vcc),
           .NS(gnd), .NZ(CI_4_6), .OP(vcc), .OS(gnd), .QC(gnd), .QR(gnd),
           .QS(gnd) );
logic2 I_51 ( .A1(vcc), .A2(gnd), .A3(A[6]), .A4(gnd), .A5(B[6]), .A6(gnd), .AZ(G6),
           .B1(gnd), .B2(gnd), .C1(B[7]), .C2(gnd), .D1(B[7]), .D2(gnd),
           .E1(vcc), .E2(gnd), .F1(vcc), .F2(gnd), .F3(A[5]), .F4(gnd),
           .F5(B[5]), .F6(gnd), .FZ(G5), .MP(gnd), .MS(A[7]), .NP(gnd),
           .NS(A[7]), .OP(vcc), .OS(gnd), .OZ(G7), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_49 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(A[4]), .A5(vcc), .A6(B[4]),
           .AZ(A4_NOR_B4), .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc),
           .D2(gnd), .E1(vcc), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(A[5]),
           .F5(vcc), .F6(B[5]), .FZ(A5_NOR_B5), .MP(vcc), .MS(gnd), .NP(vcc),
           .NS(gnd), .OP(vcc), .OS(gnd), .OZ(P5_N), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_23 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(CI), .AZ(CI0_N),
           .B1(vcc), .B2(B[0]), .C1(B[0]), .C2(gnd), .D1(B[0]), .D2(gnd),
           .E1(vcc), .E2(B[0]), .F1(vcc), .F2(gnd), .F3(vcc), .F4(gnd), .F5(gnd),
           .F6(gnd), .MP(gnd), .MS(A[0]), .NP(gnd), .NS(A[0]), .NZ(P0), .OP(vcc),
           .OS(gnd), .OZ(SUM[0]), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_21 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(G1_N), .A6(CI_2_6),
           .AZ(CI2_N), .B1(vcc), .B2(B[2]), .C1(B[2]), .C2(gnd), .D1(B[2]),
           .D2(gnd), .E1(vcc), .E2(B[2]), .F1(A[3]), .F2(gnd), .F3(B[3]),
           .F4(gnd), .F5(vcc), .F6(gnd), .FZ(A3_AND_B3), .MP(gnd), .MS(A[2]),
           .NP(gnd), .NS(A[2]), .NZ(P2), .OP(vcc), .OS(gnd), .OZ(SUM[2]),
           .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_37 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(A[2]), .A5(vcc), .A6(B[2]),
           .AZ(A2_NOR_B2), .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc),
           .D2(gnd), .E1(vcc), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(A[3]),
           .F5(vcc), .F6(B[3]), .FZ(A3_NOR_B3), .MP(vcc), .MS(gnd), .NP(vcc),
           .NS(gnd), .OP(vcc), .OS(gnd), .OZ(P3_N), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_36 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(A[0]), .A5(vcc), .A6(B[0]),
           .AZ(A0_NOR_B0), .B1(gnd), .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc),
           .D2(gnd), .E1(vcc), .E2(gnd), .F1(vcc), .F2(gnd), .F3(vcc), .F4(A[1]),
           .F5(vcc), .F6(B[1]), .FZ(A1_NOR_B1), .MP(vcc), .MS(gnd), .NP(vcc),
           .NS(gnd), .OP(vcc), .OS(gnd), .OZ(P1_N), .QC(gnd), .QR(gnd), .QS(gnd) );
logic2 I_12 ( .A1(vcc), .A2(gnd), .A3(A[2]), .A4(gnd), .A5(B[2]), .A6(gnd), .AZ(G2),
           .B1(gnd), .B2(gnd), .C1(B[3]), .C2(gnd), .D1(B[3]), .D2(gnd),
           .E1(vcc), .E2(gnd), .F1(A[3]), .F2(gnd), .F3(B[3]), .F4(gnd),
           .F5(vcc), .F6(gnd), .MP(gnd), .MS(A[3]), .NP(gnd), .NS(A[3]),
           .OP(vcc), .OS(gnd), .OZ(G3), .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // fstadd16

`endif

`ifdef fadd1_p2
`else
`define fadd1_p2
module fadd1_p2( A , B, CI, CO, S );
input A, B, CI;
output CO, S;
parameter ql_gate = `LOGIC;
supply0 GND;
supply1 VCC;

lcell2 I_6 ( .A1(GND), .A2(GND), .A3(GND), .A4(GND), .A5(GND), .A6(GND), .B1(CI),
          .B2(GND), .C1(VCC), .C2(CI), .D1(B), .D2(GND), .E1(CI), .E2(GND),
          .F1(VCC), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(B), .MP(A),
          .MS(B), .NP(A), .NS(B), .NZ(CO), .OP(GND), .OS(GND), .OZ(S), .QC(GND),
          .QR(GND), .QS(GND) );

endmodule // fadd1_p2

`endif

`ifdef ecompai
`else
`define ecompai
module ecompai( A , B, EQ2 );
 input [1:0] A;
 input [1:0] B;
output EQ2;
supply1 vcc;
supply0 gnd;

logic2 I_2 ( .A1(vcc), .A2(B[0]), .A3(vcc), .A4(gnd), .A5(vcc), .A6(gnd), .B1(gnd),
          .B2(gnd), .C1(vcc), .C2(gnd), .D1(vcc), .D2(gnd), .E1(vcc), .E2(gnd),
          .F1(vcc), .F2(B[1]), .F3(vcc), .F4(gnd), .F5(vcc), .F6(gnd), .MP(A[1]),
          .MS(B[1]), .NP(A[1]), .NS(B[1]), .OP(A[0]), .OS(B[0]), .OZ(EQ2),
          .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // ecompai

`endif

`ifdef ecompa
`else
`define ecompa
module ecompa( A , B, EQ2 );
 input [1:0] A;
 input [1:0] B;
output EQ2;
supply1 vcc;
supply0 gnd;

logic2 I_2 ( .A1(vcc), .A2(B[0]), .A3(vcc), .A4(gnd), .A5(vcc), .A6(gnd), .B1(vcc),
          .B2(gnd), .C1(gnd), .C2(gnd), .D1(gnd), .D2(gnd), .E1(gnd), .E2(gnd),
          .F1(vcc), .F2(B[1]), .F3(vcc), .F4(gnd), .F5(vcc), .F6(gnd), .MP(A[1]),
          .MS(B[1]), .NP(A[1]), .NS(B[1]), .OP(A[0]), .OS(B[0]), .OZ(EQ2),
          .QC(gnd), .QR(gnd), .QS(vcc) );

endmodule // ecompa

`endif

`ifdef ecomp8
`else
`define ecomp8
module ecomp8( A , B, EQ );
 input [7:0] A;
 input [7:0] B;
output EQ;
wire N_1;
wire N_2;
wire N_3;
wire N_4;

ecompa I_7 ( .A({ A[7:6] }), .B({ B[7:6] }), .EQ2(N_2) );
ecompa I_8 ( .A({ A[5:4] }), .B({ B[5:4] }), .EQ2(N_3) );
ecompa I_9 ( .A({ A[3:2] }), .B({ B[3:2] }), .EQ2(N_4) );
ecompa I_10 ( .A({ A[1:0] }), .B({ B[1:0] }), .EQ2(N_1) );
and4i0 I_1 ( .A(N_1), .B(N_4), .C(N_3), .D(N_2), .Q(EQ) );

endmodule // ecomp8

`endif

`ifdef ecomp4
`else
`define ecomp4
module ecomp4( A , B, EQ );
 input [3:0] A;
 input [3:0] B;
output EQ;
wire N_1;
wire N_2;

ecompa I_8 ( .A({ A[3:2] }), .B({ B[3:2] }), .EQ2(N_1) );
ecompa I_9 ( .A({ A[1:0] }), .B({ B[1:0] }), .EQ2(N_2) );
and2i0 I_7 ( .A(N_2), .B(N_1), .Q(EQ) );

endmodule // ecomp4

`endif

`ifdef ecomp32
`else
`define ecomp32
module ecomp32( A , B, EQ );
 input [31:0] A;
 input [31:0] B;
output EQ;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;
wire N_15;
wire N_16;
wire N_17;

ecompai I_35 ( .A({ A[31:30] }), .B({ B[31:30] }), .EQ2(N_17) );
ecompai I_20 ( .A({ A[29:28] }), .B({ B[29:28] }), .EQ2(N_16) );
ecompai I_21 ( .A({ A[27:26] }), .B({ B[27:26] }), .EQ2(N_15) );
ecompai I_22 ( .A({ A[25:24] }), .B({ B[25:24] }), .EQ2(N_13) );
ecompai I_23 ( .A({ A[23:22] }), .B({ B[23:22] }), .EQ2(N_11) );
ecompai I_24 ( .A({ A[21:20] }), .B({ B[21:20] }), .EQ2(N_9) );
ecompai I_19 ( .A({ A[19:18] }), .B({ B[19:18] }), .EQ2(N_7) );
ecompa I_37 ( .A({ A[17:16] }), .B({ B[17:16] }), .EQ2(N_5) );
ecompa I_36 ( .A({ A[15:14] }), .B({ B[15:14] }), .EQ2(N_2) );
ecompa I_28 ( .A({ A[13:12] }), .B({ B[13:12] }), .EQ2(N_3) );
ecompa I_34 ( .A({ A[11:10] }), .B({ B[11:10] }), .EQ2(N_4) );
ecompa I_33 ( .A({ A[9:8] }), .B({ B[9:8] }), .EQ2(N_6) );
ecompa I_32 ( .A({ A[7:6] }), .B({ B[7:6] }), .EQ2(N_8) );
ecompa I_31 ( .A({ A[5:4] }), .B({ B[5:4] }), .EQ2(N_10) );
ecompa I_30 ( .A({ A[3:2] }), .B({ B[3:2] }), .EQ2(N_12) );
ecompa I_29 ( .A({ A[1:0] }), .B({ B[1:0] }), .EQ2(N_14) );
and16i7 I_18 ( .A(N_14), .B(N_12), .C(N_10), .D(N_8), .E(N_6), .F(N_4), .G(N_3),
            .H(N_2), .I(N_5), .J(N_7), .K(N_9), .L(N_11), .M(N_13), .N(N_15),
            .O(N_16), .P(N_17), .Q(EQ) );

endmodule // ecomp32

`endif

`ifdef ecomp2
`else
`define ecomp2
module ecomp2( A , B, EQ );
 input [1:0] A;
 input [1:0] B;
output EQ;
supply1 vcc;
supply0 gnd;
wire N_1;
wire N_2;

logic2 I_3 ( .A1(A[0]), .A2(gnd), .A3(vcc), .A4(gnd), .A5(vcc), .A6(B[0]),
          .B1(B[0]), .B2(A[0]), .C1(B[0]), .C2(A[0]), .D1(vcc), .D2(A[1]),
          .E1(A[1]), .E2(gnd), .F1(vcc), .F2(gnd), .F3(N_1), .F4(gnd), .F5(vcc),
          .F6(N_2), .FZ(EQ), .MP(gnd), .MS(B[1]), .NP(gnd), .NS(B[1]), .NZ(N_1),
          .OP(vcc), .OS(gnd), .OZ(N_2), .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // ecomp2

`endif

`ifdef ecomp16
`else
`define ecomp16
module ecomp16( A , B, EQ );
 input [15:0] A;
 input [15:0] B;
output EQ;
supply1 vcc;
supply0 gnd;
wire N_66;
wire N_67;
wire N_69;
wire N_70;
wire N_72;
wire N_74;
wire N_76;
wire N_78;

ecompa I_27 ( .A({ A[15:14] }), .B({ B[15:14] }), .EQ2(N_69) );
ecompa I_21 ( .A({ A[11:10] }), .B({ B[11:10] }), .EQ2(N_70) );
ecompa I_19 ( .A({ A[13:12] }), .B({ B[13:12] }), .EQ2(N_66) );
ecompa I_22 ( .A({ A[9:8] }), .B({ B[9:8] }), .EQ2(N_72) );
ecompa I_23 ( .A({ A[7:6] }), .B({ B[7:6] }), .EQ2(N_74) );
ecompa I_24 ( .A({ A[5:4] }), .B({ B[5:4] }), .EQ2(N_76) );
ecompa I_25 ( .A({ A[3:2] }), .B({ B[3:2] }), .EQ2(N_78) );
ecompa I_26 ( .A({ A[1:0] }), .B({ B[1:0] }), .EQ2(N_67) );
and16i7 I_18 ( .A(N_67), .B(N_78), .C(N_76), .D(N_74), .E(N_72), .F(N_70), .G(N_66),
            .H(N_69), .I(vcc), .J(gnd), .K(gnd), .L(gnd), .M(gnd), .N(gnd),
            .O(gnd), .P(gnd), .Q(EQ) );

endmodule // ecomp16

`endif

`ifdef cktpadff
`else
`define cktpadff
module cktpadff( FFCLK , FFCLR, FFEN, P, FFQ, Q0, Q1, Q2 );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input FFEN;
output FFQ;
input P /* synthesis syn_isclock=1 */;
output Q0, Q1, Q2;
parameter syn_macro = 1;
parameter ql_gate = `CLOCK;

ckcell2 QL1 ( .IC(Q1), .IN(Q0), .IP(P), .IQ(FFQ), .IQC(FFCLK), .IQE(FFEN),
           .IR(FFCLR), .IZ(Q2) );

endmodule // cktpadff

`endif

`ifdef ckpadff
`else
`define ckpadff
module ckpadff( FFCLK, FFCLR, FFEN, FFQ, P, Q1 );
input FFCLK /*synthesis syn_isclock=1 */;
input FFCLR /*synthesis syn_isclock=1 */;
input FFEN;
output FFQ;
input P /*synthesis syn_isclock=1 */;
output Q1;
parameter syn_macro = 1;
parameter ql_gate = `CLOCK;

ckcell2 QL1 ( .IC(Q1), .IP(P), .IQ(FFQ), .IQC(FFCLK), .IQE(FFEN), .IR(FFCLR) );

endmodule // ckpadff

`endif

`ifdef ckdpadff
`else
`define ckdpadff
module ckdpadff( FFCLK , FFCLR, FFEN, P, FFQ, Q0, Q2 );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input FFEN;
output FFQ;
input P /* synthesis syn_isclock=1 */;
output Q0, Q2;
parameter syn_macro = 1;
parameter ql_gate = `CLOCK;

ckcell2 QL1 ( .IN(Q0), .IP(P), .IQ(FFQ), .IQC(FFCLK), .IQE(FFEN), .IR(FFCLR),
           .IZ(Q2) );

endmodule // ckdpadff

`endif

`ifdef bpad8ff
`else
`define bpad8ff
module bpad8ff( A2 , EN, FFCLK, FFCLR, FFEN, FFQ, Q, P );
 input [7:0] A2;
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input EN, FFEN;
 output [7:0] FFQ;
 inout [7:0] P;
 output [7:0] Q;

bipadff QL0 ( .A2(A2[0]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[0]), .P(P[0]), .Q(Q[0]) );
bipadff QL1 ( .A2(A2[1]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[1]), .P(P[1]), .Q(Q[1]) );
bipadff QL2 ( .A2(A2[2]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[2]), .P(P[2]), .Q(Q[2]) );
bipadff QL3 ( .A2(A2[3]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[3]), .P(P[3]), .Q(Q[3]) );
bipadff QL4 ( .A2(A2[4]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[4]), .P(P[4]), .Q(Q[4]) );
bipadff QL5 ( .A2(A2[5]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[5]), .P(P[5]), .Q(Q[5]) );
bipadff QL6 ( .A2(A2[6]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[6]), .P(P[6]), .Q(Q[6]) );
bipadff QL7 ( .A2(A2[7]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[7]), .P(P[7]), .Q(Q[7]) );

endmodule // bpad8ff

`endif

`ifdef bpad4ff
`else
`define bpad4ff
module bpad4ff( A2 , EN, FFCLK, FFCLR, FFEN, FFQ, Q, P );
 input [3:0] A2;
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input EN, FFEN;
 output [3:0] FFQ;
 inout [3:0] P;
 output [3:0] Q;

bipadff QL0 ( .A2(A2[0]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[0]), .P(P[0]), .Q(Q[0]) );
bipadff QL1 ( .A2(A2[1]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[1]), .P(P[1]), .Q(Q[1]) );
bipadff QL2 ( .A2(A2[2]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[2]), .P(P[2]), .Q(Q[2]) );
bipadff QL3 ( .A2(A2[3]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[3]), .P(P[3]), .Q(Q[3]) );

endmodule // bpad4ff

`endif

`ifdef bpad16ff
`else
`define bpad16ff
module bpad16ff( A2 , EN, FFCLK, FFCLR, FFEN, FFQ, Q, P );
 input [15:0] A2;
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input EN, FFEN;
 output [15:0] FFQ;
 inout [15:0] P;
 output [15:0] Q;

bipadff QL0 ( .A2(A2[0]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[0]), .P(P[0]), .Q(Q[0]) );
bipadff QL1 ( .A2(A2[1]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[1]), .P(P[1]), .Q(Q[1]) );
bipadff QL2 ( .A2(A2[2]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[2]), .P(P[2]), .Q(Q[2]) );
bipadff QL3 ( .A2(A2[3]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[3]), .P(P[3]), .Q(Q[3]) );
bipadff QL4 ( .A2(A2[4]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[4]), .P(P[4]), .Q(Q[4]) );
bipadff QL5 ( .A2(A2[5]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[5]), .P(P[5]), .Q(Q[5]) );
bipadff QL6 ( .A2(A2[6]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[6]), .P(P[6]), .Q(Q[6]) );
bipadff QL7 ( .A2(A2[7]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[7]), .P(P[7]), .Q(Q[7]) );
bipadff QL8 ( .A2(A2[8]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[8]), .P(P[8]), .Q(Q[8]) );
bipadff QL9 ( .A2(A2[9]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
           .FFQ(FFQ[9]), .P(P[9]), .Q(Q[9]) );
bipadff QL10 ( .A2(A2[10]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
            .FFQ(FFQ[10]), .P(P[10]), .Q(Q[10]) );
bipadff QL11 ( .A2(A2[11]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
            .FFQ(FFQ[11]), .P(P[11]), .Q(Q[11]) );
bipadff QL12 ( .A2(A2[12]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
            .FFQ(FFQ[12]), .P(P[12]), .Q(Q[12]) );
bipadff QL13 ( .A2(A2[13]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
            .FFQ(FFQ[13]), .P(P[13]), .Q(Q[13]) );
bipadff QL14 ( .A2(A2[14]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
            .FFQ(FFQ[14]), .P(P[14]), .Q(Q[14]) );
bipadff QL15 ( .A2(A2[15]), .EN(EN), .FFCLK(FFCLK), .FFCLR(FFCLR), .FFEN(FFEN),
            .FFQ(FFQ[15]), .P(P[15]), .Q(Q[15]) );

endmodule // bpad16ff

`endif

`ifdef bipadff
`else
`define bipadff
module bipadff( A2 , EN, FFCLK, FFCLR, FFEN, FFQ, Q, P );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input A2, EN, FFEN;
output FFQ;
inout P;
output Q;
parameter ql_gate = `BIDIR;
supply1 VCC;

bicell2 QL1 ( .I1(VCC), .I2(A2), .IC(FFCLK), .IE(EN), .IP(P), .IQ(FFQ), .IQE(FFEN),
           .IR(FFCLR), .IZ(Q) );

endmodule // bipadff

`endif

`ifdef biorpadf
`else
`define biorpadf
module biorpadf( A1 , A2, EN, FFCLK, FFCLR, FFEN, FFQ, Q, P );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input A1, A2, EN, FFEN;
output FFQ;
inout P;
output Q;
parameter ql_gate = `BIDIR;

bicell2 QL1 ( .I1(A1), .I2(A2), .IC(FFCLK), .IE(EN), .IP(P), .IQ(FFQ), .IQE(FFEN),
           .IR(FFCLR), .IZ(Q) );

endmodule // biorpadf

`endif

`ifdef biipadff
`else
`define biipadff
module biipadff( A1 , EN, FFCLK, FFCLR, FFEN, FFQ, Q, P );
input FFCLK /* synthesis syn_isclock=1 */;
input FFCLR /* synthesis syn_isclock=1 */;
input A1, EN, FFEN;
output FFQ;
inout P;
output Q;
parameter ql_gate = `BIDIR;
supply0 gnd;

bicell2 QL1 ( .I1(A1), .I2(gnd), .IC(FFCLK), .IE(EN), .IP(P), .IQ(FFQ), .IQE(FFEN),
           .IR(FFCLR), .IZ(Q) );

endmodule // biipadff

`endif

`ifdef and9i4
`else
`define and9i4
module and9i4( A , B, C, D, E, F, G, H, I, Q );
input A, B, C, D, E, F, G, H, I;
output Q;
supply0 GND;
supply1 VCC;

logic2 I_1 ( .A1(GND), .A2(GND), .A3(GND), .A4(GND), .A5(GND), .A6(GND), .B1(GND),
          .B2(GND), .C1(GND), .C2(GND), .D1(GND), .D2(GND), .E1(A), .E2(F),
          .F1(C), .F2(G), .F3(D), .F4(H), .F5(E), .F6(I), .MP(GND), .MS(GND),
          .NP(B), .NS(GND), .NZ(Q), .OP(VCC), .OS(GND), .QC(GND), .QR(GND),
          .QS(GND) );

endmodule // and9i4

`endif

`ifdef and8i1
`else
`define and8i1
module and8i1( A , B, C, D, E, F, G, H, Q );
input A, B, C, D, E, F, G, H;
output Q;
supply0 GND;
supply1 VCC;

logic2 I_1 ( .A1(VCC), .A2(A), .A3(B), .A4(GND), .A5(C), .A6(GND), .B1(GND),
          .B2(GND), .C1(GND), .C2(GND), .D1(GND), .D2(GND), .E1(VCC), .E2(GND),
          .F1(F), .F2(GND), .F3(G), .F4(GND), .F5(H), .F6(GND), .MP(GND),
          .MS(GND), .NP(E), .NS(GND), .OP(D), .OS(GND), .OZ(Q), .QC(GND),
          .QR(GND), .QS(GND) );

endmodule // and8i1

`endif

`ifdef and8i0
`else
`define and8i0
module and8i0( A , B, C, D, E, F, G, H, Q );
input A, B, C, D, E, F, G, H;
output Q;
supply0 GND;
supply1 VCC;

logic2 I_1 ( .A1(A), .A2(GND), .A3(B), .A4(GND), .A5(C), .A6(GND), .B1(GND),
          .B2(GND), .C1(GND), .C2(GND), .D1(GND), .D2(GND), .E1(VCC), .E2(GND),
          .F1(F), .F2(GND), .F3(G), .F4(GND), .F5(H), .F6(GND), .MP(GND),
          .MS(GND), .NP(E), .NS(GND), .OP(D), .OS(GND), .OZ(Q), .QC(GND),
          .QR(GND), .QS(GND) );

endmodule // and8i0

`endif

`ifdef and7i1
`else
`define and7i1
module and7i1( A , B, C, D, E, F, G, Q );
input A, B, C, D, E, F, G;
output Q;
supply0 GND;
supply1 VCC;

logic2 I_1 ( .A1(A), .A2(GND), .A3(B), .A4(GND), .A5(C), .A6(GND), .B1(GND),
          .B2(GND), .C1(GND), .C2(GND), .D1(GND), .D2(GND), .E1(VCC), .E2(GND),
          .F1(F), .F2(GND), .F3(VCC), .F4(G), .F5(D), .F6(GND), .MP(GND),
          .MS(GND), .NP(E), .NS(GND), .OP(VCC), .OS(GND), .OZ(Q), .QC(GND),
          .QR(GND), .QS(GND) );

endmodule // and7i1

`endif

`ifdef and7i0
`else
`define and7i0
module and7i0( A , B, C, D, E, F, G, Q );
input A, B, C, D, E, F, G;
output Q;
supply0 GND;
supply1 VCC;

logic2 I_1 ( .A1(A), .A2(GND), .A3(B), .A4(GND), .A5(C), .A6(GND), .B1(GND),
          .B2(GND), .C1(GND), .C2(GND), .D1(GND), .D2(GND), .E1(VCC), .E2(GND),
          .F1(F), .F2(GND), .F3(G), .F4(GND), .F5(D), .F6(GND), .MP(GND),
          .MS(GND), .NP(E), .NS(GND), .OP(VCC), .OS(GND), .OZ(Q), .QC(GND),
          .QR(GND), .QS(GND) );

endmodule // and7i0

`endif

`ifdef and16i7
`else
`define and16i7
module and16i7( A , B, C, D, E, F, G, H, I, J, K, L, M, N, O, P, Q );
input A, B, C, D, E, F, G, H, I, J, K, L, M, N, O, P;
output Q;
supply0 gnd;

logic2 I_3 ( .A1(A), .A2(J), .A3(B), .A4(K), .A5(C), .A6(L), .B1(gnd), .B2(gnd),
          .C1(gnd), .C2(gnd), .D1(gnd), .D2(gnd), .E1(E), .E2(M), .F1(G), .F2(N),
          .F3(H), .F4(O), .F5(I), .F6(P), .MP(gnd), .MS(gnd), .NP(F), .NS(gnd),
          .OP(D), .OS(gnd), .OZ(Q), .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // and16i7

`endif

`ifdef shft8
`else
`define shft8
module shft8( CLK , CLR, D, EN, LOAD, SI, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [7:0] D;
input EN, LOAD;
 output [7:0] Q;
input SI;

shft4 QL2 ( .CLK(CLK), .CLR(CLR), .D({ D[7:4] }), .EN(EN), .LOAD(LOAD),
         .Q({ Q[7:4] }), .SI(Q[3]) );
shft4 QL1 ( .CLK(CLK), .CLR(CLR), .D({ D[3:0] }), .EN(EN), .LOAD(LOAD),
         .Q({ Q[3:0] }), .SI(SI) );

endmodule // shft8

`endif

`ifdef shft4
`else
`define shft4
module shft4( CLK , CLR, D, EN, LOAD, SI, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [3:0] D;
input EN, LOAD;
 output [3:0] Q;
input SI;

shiftbit QL1 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .EN(EN), .LOAD(LOAD), .Q(Q[0]),
            .SI(SI) );
shiftbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .EN(EN), .LOAD(LOAD), .Q(Q[1]),
            .SI(Q[0]) );
shiftbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .EN(EN), .LOAD(LOAD), .Q(Q[2]),
            .SI(Q[1]) );
shiftbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .EN(EN), .LOAD(LOAD), .Q(Q[3]),
            .SI(Q[2]) );

endmodule // shft4

`endif

`ifdef shft16
`else
`define shft16
module shft16( CLK , CLR, D, EN, LOAD, SI, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [15:0] D;
input EN, LOAD;
 output [15:0] Q;
input SI;

shft4 QL4 ( .CLK(CLK), .CLR(CLR), .D({ D[15:12] }), .EN(EN), .LOAD(LOAD),
         .Q({ Q[15:12] }), .SI(Q[11]) );
shft4 QL3 ( .CLK(CLK), .CLR(CLR), .D({ D[11:8] }), .EN(EN), .LOAD(LOAD),
         .Q({ Q[11:8] }), .SI(Q[7]) );
shft4 QL2 ( .CLK(CLK), .CLR(CLR), .D({ D[7:4] }), .EN(EN), .LOAD(LOAD),
         .Q({ Q[7:4] }), .SI(Q[3]) );
shft4 QL1 ( .CLK(CLK), .CLR(CLR), .D({ D[3:0] }), .EN(EN), .LOAD(LOAD),
         .Q({ Q[3:0] }), .SI(SI) );

endmodule // shft16

`endif

`ifdef bshft8
`else
`define bshft8
module bshft8( CLK , CLR, D, LSI, RSI, S0, S1, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [7:0] D;
input LSI;
 output [7:0] Q;
input RSI, S0, S1;

bshft4 QL2 ( .CLK(CLK), .CLR(CLR), .D({ D[7:4] }), .LSI(Q[3]), .Q({ Q[7:4] }),
          .RSI(RSI), .S0(S0), .S1(S1) );
bshft4 QL1 ( .CLK(CLK), .CLR(CLR), .D({ D[3:0] }), .LSI(LSI), .Q({ Q[3:0] }),
          .RSI(Q[4]), .S0(S0), .S1(S1) );

endmodule // bshft8

`endif

`ifdef bshft4
`else
`define bshft4
module bshft4( CLK , CLR, D, LSI, RSI, S0, S1, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [3:0] D;
input LSI;
 output [3:0] Q;
input RSI, S0, S1;

bishbit QL1 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .LSI(LSI), .Q(Q[0]), .RSI(Q[1]),
           .S0(S0), .S1(S1) );
bishbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .LSI(Q[1]), .Q(Q[2]), .RSI(Q[3]),
           .S0(S0), .S1(S1) );
bishbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .LSI(Q[0]), .Q(Q[1]), .RSI(Q[2]),
           .S0(S0), .S1(S1) );
bishbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .LSI(Q[2]), .Q(Q[3]), .RSI(RSI),
           .S0(S0), .S1(S1) );

endmodule // bshft4

`endif

`ifdef bshft16
`else
`define bshft16
module bshft16( CLK , CLR, D, LSI, RSI, S0, S1, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [15:0] D;
input LSI;
 output [15:0] Q;
input RSI, S0, S1;

bshft4 QL4 ( .CLK(CLK), .CLR(CLR), .D({ D[15:12] }), .LSI(Q[11]),
          .Q({ Q[15:12] }), .RSI(RSI), .S0(S0), .S1(S1) );
bshft4 QL3 ( .CLK(CLK), .CLR(CLR), .D({ D[11:8] }), .LSI(Q[7]), .Q({ Q[11:8] }),
          .RSI(Q[12]), .S0(S0), .S1(S1) );
bshft4 QL2 ( .CLK(CLK), .CLR(CLR), .D({ D[7:4] }), .LSI(Q[3]), .Q({ Q[7:4] }),
          .RSI(Q[8]), .S0(S0), .S1(S1) );
bshft4 QL1 ( .CLK(CLK), .CLR(CLR), .D({ D[3:0] }), .LSI(LSI), .Q({ Q[3:0] }),
          .RSI(Q[4]), .S0(S0), .S1(S1) );

endmodule // bshft16

`endif

`ifdef rgec8
`else
`define rgec8
module rgec8( CLK , CLR, D, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [7:0] D;
input EN;
 output [7:0] Q;
supply0 GND;

dffepc QL8 ( .CLK(CLK), .CLR(CLR), .D(D[4]), .EN(EN), .PRE(GND), .Q(Q[4]) );
dffepc QL7 ( .CLK(CLK), .CLR(CLR), .D(D[5]), .EN(EN), .PRE(GND), .Q(Q[5]) );
dffepc QL6 ( .CLK(CLK), .CLR(CLR), .D(D[6]), .EN(EN), .PRE(GND), .Q(Q[6]) );
dffepc QL5 ( .CLK(CLK), .CLR(CLR), .D(D[7]), .EN(EN), .PRE(GND), .Q(Q[7]) );
dffepc QL4 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .EN(EN), .PRE(GND), .Q(Q[0]) );
dffepc QL3 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .EN(EN), .PRE(GND), .Q(Q[1]) );
dffepc QL2 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .EN(EN), .PRE(GND), .Q(Q[2]) );
dffepc QL1 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .EN(EN), .PRE(GND), .Q(Q[3]) );

endmodule // rgec8

`endif

`ifdef rgec4
`else
`define rgec4
module rgec4( CLK , CLR, D, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [3:0] D;
input EN;
 output [3:0] Q;
supply0 GND;

dffepc QL4 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .EN(EN), .PRE(GND), .Q(Q[0]) );
dffepc QL3 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .EN(EN), .PRE(GND), .Q(Q[1]) );
dffepc QL2 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .EN(EN), .PRE(GND), .Q(Q[2]) );
dffepc QL1 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .EN(EN), .PRE(GND), .Q(Q[3]) );

endmodule // rgec4

`endif

`ifdef rgec16
`else
`define rgec16
module rgec16( CLK , CLR, D, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [15:0] D;
input EN;
 output [15:0] Q;
supply0 GND;

dffepc QL16 ( .CLK(CLK), .CLR(CLR), .D(D[12]), .EN(EN), .PRE(GND), .Q(Q[12]) );
dffepc QL15 ( .CLK(CLK), .CLR(CLR), .D(D[13]), .EN(EN), .PRE(GND), .Q(Q[13]) );
dffepc QL14 ( .CLK(CLK), .CLR(CLR), .D(D[14]), .EN(EN), .PRE(GND), .Q(Q[14]) );
dffepc QL13 ( .CLK(CLK), .CLR(CLR), .D(D[15]), .EN(EN), .PRE(GND), .Q(Q[15]) );
dffepc QL12 ( .CLK(CLK), .CLR(CLR), .D(D[8]), .EN(EN), .PRE(GND), .Q(Q[8]) );
dffepc QL11 ( .CLK(CLK), .CLR(CLR), .D(D[9]), .EN(EN), .PRE(GND), .Q(Q[9]) );
dffepc QL10 ( .CLK(CLK), .CLR(CLR), .D(D[10]), .EN(EN), .PRE(GND), .Q(Q[10]) );
dffepc QL9 ( .CLK(CLK), .CLR(CLR), .D(D[11]), .EN(EN), .PRE(GND), .Q(Q[11]) );
dffepc QL8 ( .CLK(CLK), .CLR(CLR), .D(D[4]), .EN(EN), .PRE(GND), .Q(Q[4]) );
dffepc QL7 ( .CLK(CLK), .CLR(CLR), .D(D[5]), .EN(EN), .PRE(GND), .Q(Q[5]) );
dffepc QL6 ( .CLK(CLK), .CLR(CLR), .D(D[6]), .EN(EN), .PRE(GND), .Q(Q[6]) );
dffepc QL5 ( .CLK(CLK), .CLR(CLR), .D(D[7]), .EN(EN), .PRE(GND), .Q(Q[7]) );
dffepc QL4 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .EN(EN), .PRE(GND), .Q(Q[0]) );
dffepc QL3 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .EN(EN), .PRE(GND), .Q(Q[1]) );
dffepc QL2 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .EN(EN), .PRE(GND), .Q(Q[2]) );
dffepc QL1 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .EN(EN), .PRE(GND), .Q(Q[3]) );

endmodule // rgec16

`endif

`ifdef rge8
`else
`define rge8
module rge8( CLK , D, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
 input [7:0] D;
input EN;
 output [7:0] Q;

dffe QL8 ( .CLK(CLK), .D(D[0]), .EN(EN), .Q(Q[0]) );
dffe QL7 ( .CLK(CLK), .D(D[1]), .EN(EN), .Q(Q[1]) );
dffe QL6 ( .CLK(CLK), .D(D[2]), .EN(EN), .Q(Q[2]) );
dffe QL5 ( .CLK(CLK), .D(D[3]), .EN(EN), .Q(Q[3]) );
dffe QL4 ( .CLK(CLK), .D(D[4]), .EN(EN), .Q(Q[4]) );
dffe QL3 ( .CLK(CLK), .D(D[5]), .EN(EN), .Q(Q[5]) );
dffe QL2 ( .CLK(CLK), .D(D[6]), .EN(EN), .Q(Q[6]) );
dffe QL1 ( .CLK(CLK), .D(D[7]), .EN(EN), .Q(Q[7]) );

endmodule // rge8

`endif

`ifdef rge4
`else
`define rge4
module rge4( CLK , D, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
 input [3:0] D;
input EN;
 output [3:0] Q;

dffe QL1 ( .CLK(CLK), .D(D[3]), .EN(EN), .Q(Q[3]) );
dffe QL2 ( .CLK(CLK), .D(D[2]), .EN(EN), .Q(Q[2]) );
dffe QL3 ( .CLK(CLK), .D(D[1]), .EN(EN), .Q(Q[1]) );
dffe QL4 ( .CLK(CLK), .D(D[0]), .EN(EN), .Q(Q[0]) );

endmodule // rge4

`endif

`ifdef rge16
`else
`define rge16
module rge16( CLK , D, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
 input [15:0] D;
input EN;
 output [15:0] Q;

dffe QL16 ( .CLK(CLK), .D(D[0]), .EN(EN), .Q(Q[0]) );
dffe QL15 ( .CLK(CLK), .D(D[1]), .EN(EN), .Q(Q[1]) );
dffe QL14 ( .CLK(CLK), .D(D[2]), .EN(EN), .Q(Q[2]) );
dffe QL13 ( .CLK(CLK), .D(D[3]), .EN(EN), .Q(Q[3]) );
dffe QL12 ( .CLK(CLK), .D(D[4]), .EN(EN), .Q(Q[4]) );
dffe QL11 ( .CLK(CLK), .D(D[5]), .EN(EN), .Q(Q[5]) );
dffe QL10 ( .CLK(CLK), .D(D[6]), .EN(EN), .Q(Q[6]) );
dffe QL9 ( .CLK(CLK), .D(D[7]), .EN(EN), .Q(Q[7]) );
dffe QL8 ( .CLK(CLK), .D(D[8]), .EN(EN), .Q(Q[8]) );
dffe QL7 ( .CLK(CLK), .D(D[9]), .EN(EN), .Q(Q[9]) );
dffe QL6 ( .CLK(CLK), .D(D[10]), .EN(EN), .Q(Q[10]) );
dffe QL5 ( .CLK(CLK), .D(D[11]), .EN(EN), .Q(Q[11]) );
dffe QL4 ( .CLK(CLK), .D(D[12]), .EN(EN), .Q(Q[12]) );
dffe QL3 ( .CLK(CLK), .D(D[13]), .EN(EN), .Q(Q[13]) );
dffe QL2 ( .CLK(CLK), .D(D[14]), .EN(EN), .Q(Q[14]) );
dffe QL1 ( .CLK(CLK), .D(D[15]), .EN(EN), .Q(Q[15]) );

endmodule // rge16

`endif

`ifdef rgc8
`else
`define rgc8
module rgc8( CLK , CLR, D, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [7:0] D;
 output [7:0] Q;

dffc QL8 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .Q(Q[0]) );
dffc QL7 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .Q(Q[1]) );
dffc QL6 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .Q(Q[2]) );
dffc QL5 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .Q(Q[3]) );
dffc QL4 ( .CLK(CLK), .CLR(CLR), .D(D[4]), .Q(Q[4]) );
dffc QL3 ( .CLK(CLK), .CLR(CLR), .D(D[5]), .Q(Q[5]) );
dffc QL2 ( .CLK(CLK), .CLR(CLR), .D(D[6]), .Q(Q[6]) );
dffc QL1 ( .CLK(CLK), .CLR(CLR), .D(D[7]), .Q(Q[7]) );

endmodule // rgc8

`endif

`ifdef rgc4
`else
`define rgc4
module rgc4( CLK , CLR, D, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [3:0] D;
 output [3:0] Q;

dffc QL4 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .Q(Q[0]) );
dffc QL3 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .Q(Q[1]) );
dffc QL2 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .Q(Q[2]) );
dffc QL1 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .Q(Q[3]) );

endmodule // rgc4

`endif

`ifdef rgc16
`else
`define rgc16
module rgc16( CLK , CLR, D, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [15:0] D;
 output [15:0] Q;

dffc QL16 ( .CLK(CLK), .CLR(CLR), .D(D[15]), .Q(Q[15]) );
dffc QL15 ( .CLK(CLK), .CLR(CLR), .D(D[14]), .Q(Q[14]) );
dffc QL14 ( .CLK(CLK), .CLR(CLR), .D(D[13]), .Q(Q[13]) );
dffc QL13 ( .CLK(CLK), .CLR(CLR), .D(D[12]), .Q(Q[12]) );
dffc QL12 ( .CLK(CLK), .CLR(CLR), .D(D[11]), .Q(Q[11]) );
dffc QL11 ( .CLK(CLK), .CLR(CLR), .D(D[10]), .Q(Q[10]) );
dffc QL10 ( .CLK(CLK), .CLR(CLR), .D(D[9]), .Q(Q[9]) );
dffc QL9 ( .CLK(CLK), .CLR(CLR), .D(D[8]), .Q(Q[8]) );
dffc QL8 ( .CLK(CLK), .CLR(CLR), .D(D[7]), .Q(Q[7]) );
dffc QL7 ( .CLK(CLK), .CLR(CLR), .D(D[6]), .Q(Q[6]) );
dffc QL6 ( .CLK(CLK), .CLR(CLR), .D(D[5]), .Q(Q[5]) );
dffc QL5 ( .CLK(CLK), .CLR(CLR), .D(D[4]), .Q(Q[4]) );
dffc QL4 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .Q(Q[3]) );
dffc QL3 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .Q(Q[2]) );
dffc QL2 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .Q(Q[1]) );
dffc QL1 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .Q(Q[0]) );

endmodule // rgc16

`endif

`ifdef rg8
`else
`define rg8
module rg8( CLK , D, Q );
input CLK /* synthesis syn_isclock=1 */;
 input [7:0] D;
 output [7:0] Q;

dff QL7 ( .CLK(CLK), .D(D[0]), .Q(Q[0]) );
dff QL6 ( .CLK(CLK), .D(D[1]), .Q(Q[1]) );
dff QL5 ( .CLK(CLK), .D(D[2]), .Q(Q[2]) );
dff QL4 ( .CLK(CLK), .D(D[3]), .Q(Q[3]) );
dff QL3 ( .CLK(CLK), .D(D[4]), .Q(Q[4]) );
dff QL2 ( .CLK(CLK), .D(D[5]), .Q(Q[5]) );
dff QL1 ( .CLK(CLK), .D(D[6]), .Q(Q[6]) );
dff QL8 ( .CLK(CLK), .D(D[7]), .Q(Q[7]) );

endmodule // rg8

`endif

`ifdef rg4
`else
`define rg4
module rg4( CLK , D, Q );
input CLK /* synthesis syn_isclock=1 */;
 input [3:0] D;
 output [3:0] Q;

dff QL4 ( .CLK(CLK), .D(D[0]), .Q(Q[0]) );
dff QL3 ( .CLK(CLK), .D(D[1]), .Q(Q[1]) );
dff QL2 ( .CLK(CLK), .D(D[2]), .Q(Q[2]) );
dff QL1 ( .CLK(CLK), .D(D[3]), .Q(Q[3]) );

endmodule // rg4

`endif

`ifdef rg16
`else
`define rg16
module rg16( CLK , D, Q );
input CLK /* synthesis syn_isclock=1 */;
 input [15:0] D;
 output [15:0] Q;

dff QL16 ( .CLK(CLK), .D(D[0]), .Q(Q[0]) );
dff QL15 ( .CLK(CLK), .D(D[1]), .Q(Q[1]) );
dff QL14 ( .CLK(CLK), .D(D[2]), .Q(Q[2]) );
dff QL13 ( .CLK(CLK), .D(D[3]), .Q(Q[3]) );
dff QL12 ( .CLK(CLK), .D(D[4]), .Q(Q[4]) );
dff QL11 ( .CLK(CLK), .D(D[5]), .Q(Q[5]) );
dff QL10 ( .CLK(CLK), .D(D[6]), .Q(Q[6]) );
dff QL9 ( .CLK(CLK), .D(D[7]), .Q(Q[7]) );
dff QL8 ( .CLK(CLK), .D(D[8]), .Q(Q[8]) );
dff QL7 ( .CLK(CLK), .D(D[9]), .Q(Q[9]) );
dff QL6 ( .CLK(CLK), .D(D[10]), .Q(Q[10]) );
dff QL5 ( .CLK(CLK), .D(D[11]), .Q(Q[11]) );
dff QL4 ( .CLK(CLK), .D(D[12]), .Q(Q[12]) );
dff QL3 ( .CLK(CLK), .D(D[13]), .Q(Q[13]) );
dff QL2 ( .CLK(CLK), .D(D[14]), .Q(Q[14]) );
dff QL1 ( .CLK(CLK), .D(D[15]), .Q(Q[15]) );

endmodule // rg16

`endif

`ifdef tripados
`else
`define tripados
module tripados( EN , P );
input EN;
output P;
parameter ql_gate = `BIDIR;
supply1 VCC;
supply0 GND;

bicell QL1 ( .I1(GND), .I2(VCC), .IE(EN), .IP(P) );

endmodule // tripados

`endif

`ifdef tripadod
`else
`define tripadod
module tripadod( EN , P );
input EN;
output P;
parameter ql_gate = `BIDIR;
supply1 VCC;
supply0 GND;

bicell QL1 ( .I1(VCC), .I2(GND), .IE(EN), .IP(P) );

endmodule // tripadod

`endif

`ifdef tripad
`else
`define tripad
module tripad( A , EN, P );
input A, EN;
output P;
parameter ql_gate = `BIDIR;
supply1 VCC;

bicell QL1 ( .I1(VCC), .I2(A), .IE(EN), .IP(P) );

endmodule // tripad

`endif

`ifdef triorpad
`else
`define triorpad
module triorpad( A1 , A2, EN, P );
input A1, A2, EN;
output P;
parameter ql_gate = `BIDIR;

bicell QL1 ( .I1(A1), .I2(A2), .IE(EN), .IP(P) );

endmodule // triorpad

`endif

`ifdef triipad
`else
`define triipad
module triipad( A , EN, P );
input A, EN;
output P;
parameter ql_gate = `BIDIR;
supply0 GND;

bicell QL1 ( .I1(A), .I2(GND), .IE(EN), .IP(P) );

endmodule // triipad

`endif

`ifdef tpad8
`else
`define tpad8
module tpad8( A , EN, P );
 input [7:0] A;
input EN;
 output [7:0] P;

tripad QL1 ( .A(A[0]), .EN(EN), .P(P[0]) );
tripad QL2 ( .A(A[1]), .EN(EN), .P(P[1]) );
tripad QL3 ( .A(A[2]), .EN(EN), .P(P[2]) );
tripad QL4 ( .A(A[3]), .EN(EN), .P(P[3]) );
tripad QL5 ( .A(A[4]), .EN(EN), .P(P[4]) );
tripad QL6 ( .A(A[5]), .EN(EN), .P(P[5]) );
tripad QL7 ( .A(A[6]), .EN(EN), .P(P[6]) );
tripad QL8 ( .A(A[7]), .EN(EN), .P(P[7]) );

endmodule // tpad8

`endif

`ifdef tpad4
`else
`define tpad4
module tpad4( A , EN, P );
 input [3:0] A;
input EN;
 output [3:0] P;

tripad QL1 ( .A(A[0]), .EN(EN), .P(P[0]) );
tripad QL2 ( .A(A[1]), .EN(EN), .P(P[1]) );
tripad QL3 ( .A(A[2]), .EN(EN), .P(P[2]) );
tripad QL4 ( .A(A[3]), .EN(EN), .P(P[3]) );

endmodule // tpad4

`endif

`ifdef tpad16
`else
`define tpad16
module tpad16( A , EN, P );
 input [15:0] A;
input EN;
 output [15:0] P;

tripad QL1 ( .A(A[15]), .EN(EN), .P(P[15]) );
tripad QL2 ( .A(A[14]), .EN(EN), .P(P[14]) );
tripad QL3 ( .A(A[13]), .EN(EN), .P(P[13]) );
tripad QL4 ( .A(A[12]), .EN(EN), .P(P[12]) );
tripad QL5 ( .A(A[11]), .EN(EN), .P(P[11]) );
tripad QL6 ( .A(A[10]), .EN(EN), .P(P[10]) );
tripad QL7 ( .A(A[9]), .EN(EN), .P(P[9]) );
tripad QL8 ( .A(A[8]), .EN(EN), .P(P[8]) );
tripad QL9 ( .A(A[7]), .EN(EN), .P(P[7]) );
tripad QL10 ( .A(A[6]), .EN(EN), .P(P[6]) );
tripad QL11 ( .A(A[5]), .EN(EN), .P(P[5]) );
tripad QL12 ( .A(A[4]), .EN(EN), .P(P[4]) );
tripad QL13 ( .A(A[3]), .EN(EN), .P(P[3]) );
tripad QL14 ( .A(A[2]), .EN(EN), .P(P[2]) );
tripad QL15 ( .A(A[1]), .EN(EN), .P(P[1]) );
tripad QL16 ( .A(A[0]), .EN(EN), .P(P[0]) );

endmodule // tpad16

`endif

`ifdef outpad
`else
`define outpad
module outpad( A , P );
input A;
output P;
parameter ql_gate = `BIDIR;
supply1 VCC;

bicell QL1 ( .I1(VCC), .I2(A), .IE(VCC), .IP(P) );

endmodule // outpad

`endif

`ifdef outorpad
`else
`define outorpad
module outorpad( A1 , A2, P );
input A1, A2;
output P;
parameter ql_gate = `BIDIR;
supply1 VCC;

bicell QL1 ( .I1(A1), .I2(A2), .IE(VCC), .IP(P) );

endmodule // outorpad

`endif

`ifdef outipad
`else
`define outipad
module outipad( A , P );
input A;
output P;
parameter ql_gate = `BIDIR;
supply1 VCC;
supply0 GND;

bicell QL1 ( .I1(A), .I2(GND), .IE(VCC), .IP(P) );

endmodule // outipad

`endif

`ifdef opad8
`else
`define opad8
module opad8( A , P );
 input [7:0] A;
 output [7:0] P;

outpad QL1 ( .A(A[3]), .P(P[3]) );
outpad QL2 ( .A(A[2]), .P(P[2]) );
outpad QL3 ( .A(A[1]), .P(P[1]) );
outpad QL4 ( .A(A[0]), .P(P[0]) );
outpad QL5 ( .A(A[7]), .P(P[7]) );
outpad QL6 ( .A(A[6]), .P(P[6]) );
outpad QL7 ( .A(A[5]), .P(P[5]) );
outpad QL8 ( .A(A[4]), .P(P[4]) );

endmodule // opad8

`endif

`ifdef opad4
`else
`define opad4
module opad4( A , P );
 input [3:0] A;
 output [3:0] P;

outpad QL1 ( .A(A[3]), .P(P[3]) );
outpad QL2 ( .A(A[2]), .P(P[2]) );
outpad QL3 ( .A(A[1]), .P(P[1]) );
outpad QL4 ( .A(A[0]), .P(P[0]) );

endmodule // opad4

`endif

`ifdef opad16
`else
`define opad16
module opad16( A , P );
 input [15:0] A;
 output [15:0] P;

outpad QL1 ( .A(A[15]), .P(P[15]) );
outpad QL2 ( .A(A[12]), .P(P[12]) );
outpad QL3 ( .A(A[13]), .P(P[13]) );
outpad QL4 ( .A(A[14]), .P(P[14]) );
outpad QL5 ( .A(A[11]), .P(P[11]) );
outpad QL6 ( .A(A[10]), .P(P[10]) );
outpad QL7 ( .A(A[9]), .P(P[9]) );
outpad QL8 ( .A(A[8]), .P(P[8]) );
outpad QL9 ( .A(A[4]), .P(P[4]) );
outpad QL10 ( .A(A[5]), .P(P[5]) );
outpad QL11 ( .A(A[6]), .P(P[6]) );
outpad QL12 ( .A(A[7]), .P(P[7]) );
outpad QL13 ( .A(A[0]), .P(P[0]) );
outpad QL14 ( .A(A[1]), .P(P[1]) );
outpad QL15 ( .A(A[2]), .P(P[2]) );
outpad QL16 ( .A(A[3]), .P(P[3]) );

endmodule // opad16

`endif

`ifdef ipad8
`else
`define ipad8
module ipad8( P , Q );
 input [7:0] P;
 output [7:0] Q;

inpad QL1 ( .P(P[3]), .Q(Q[3]) );
inpad QL2 ( .P(P[2]), .Q(Q[2]) );
inpad QL3 ( .P(P[1]), .Q(Q[1]) );
inpad QL4 ( .P(P[0]), .Q(Q[0]) );
inpad QL5 ( .P(P[7]), .Q(Q[7]) );
inpad QL6 ( .P(P[6]), .Q(Q[6]) );
inpad QL7 ( .P(P[5]), .Q(Q[5]) );
inpad QL8 ( .P(P[4]), .Q(Q[4]) );

endmodule // ipad8

`endif

`ifdef ipad4
`else
`define ipad4
module ipad4( P , Q );
 input [3:0] P;
 output [3:0] Q;

inpad QL1 ( .P(P[3]), .Q(Q[3]) );
inpad QL2 ( .P(P[2]), .Q(Q[2]) );
inpad QL3 ( .P(P[1]), .Q(Q[1]) );
inpad QL4 ( .P(P[0]), .Q(Q[0]) );

endmodule // ipad4

`endif

`ifdef ipad16
`else
`define ipad16
module ipad16( P , Q );
 input [15:0] P;
 output [15:0] Q;

inpad QL1 ( .P(P[15]), .Q(Q[15]) );
inpad QL2 ( .P(P[12]), .Q(Q[12]) );
inpad QL3 ( .P(P[13]), .Q(Q[13]) );
inpad QL4 ( .P(P[14]), .Q(Q[14]) );
inpad QL5 ( .P(P[11]), .Q(Q[11]) );
inpad QL6 ( .P(P[10]), .Q(Q[10]) );
inpad QL7 ( .P(P[9]), .Q(Q[9]) );
inpad QL8 ( .P(P[8]), .Q(Q[8]) );
inpad QL9 ( .P(P[4]), .Q(Q[4]) );
inpad QL10 ( .P(P[5]), .Q(Q[5]) );
inpad QL11 ( .P(P[6]), .Q(Q[6]) );
inpad QL12 ( .P(P[7]), .Q(Q[7]) );
inpad QL13 ( .P(P[0]), .Q(Q[0]) );
inpad QL14 ( .P(P[1]), .Q(Q[1]) );
inpad QL15 ( .P(P[2]), .Q(Q[2]) );
inpad QL16 ( .P(P[3]), .Q(Q[3]) );

endmodule // ipad16

`endif

`ifdef inpad
`else
`define inpad
module inpad( P , Q );
input P;
output Q;
parameter ql_gate = `BIDIR;
supply1 VCC;
supply0 GND;

bicell QL1 ( .I1(GND), .I2(VCC), .IE(GND), .IP(P), .IZ(Q) );

endmodule // inpad

`endif

`ifdef hdpad
`else
`define hdpad
module hdpad( P , Q );
input P;
output Q;
parameter syn_macro = 1;
parameter ql_gate = `INCELL;

incell QL1 ( .IP(P), .IZ(Q) );

endmodule // hdpad

`endif

`ifdef hdipad
`else
`define hdipad
module hdipad( P , Q );
input P;
output Q;
parameter ql_gate = `INCELL;

incell QL1 ( .IN(Q), .IP(P) );

endmodule // hdipad

`endif

`ifdef hddpad
`else
`define hddpad
module hddpad( P , Q0, Q1 );
input P;
output Q0, Q1;
parameter syn_macro = 1;
parameter ql_gate = `INCELL;

incell QL1 ( .IN(Q0), .IP(P), .IZ(Q1) );

endmodule // hddpad

`endif

`ifdef hd3pad
`else
`define hd3pad
module hd3pad( P , Q ) /* synthesis syn_black_box black_box_tri_pins="Q" */;
input P;
output Q;
parameter syn_macro = 1;

hdpad QL1 ( .P(P), .Q(Q) );
hdpad QL2 ( .P(P), .Q(Q) );
hdpad QL3 ( .P(P), .Q(Q) );

endmodule // hd3pad

`endif

`ifdef hd2pad
`else
`define hd2pad
module hd2pad( P , Q ) /* synthesis syn_black_box black_box_tri_pins="Q" */;
input P;
output Q;
parameter syn_macro = 1;

hdpad QL1 ( .P(P), .Q(Q) );
hdpad QL2 ( .P(P), .Q(Q) );

endmodule // hd2pad

`endif

`ifdef cktpad
`else
`define cktpad
module cktpad( P , Q0, Q1, Q2 );
input P /*synthesis syn_isclock=1 */;
output Q0, Q1, Q2;
parameter syn_macro = 1;
parameter ql_gate = `CLOCK;

ckcell QL1 ( .IC(Q1), .IN(Q0), .IP(P), .IZ(Q2) );

endmodule // cktpad

`endif

`ifdef ckpad
`else
`define ckpad
module ckpad( P , Q );
input P /*synthesis syn_isclock=1 */;
output Q;
parameter ql_gate = `CLOCK;

ckcell QL1 ( .IC(Q), .IP(P) );

endmodule // ckpad

`endif

`ifdef ckdpad
`else
`define ckdpad
module ckdpad( P , Q0, Q2 );
input P /*synthesis syn_isclock=1 */;
output Q0, Q2;
parameter syn_macro = 1;
parameter ql_gate = `CLOCK;

ckcell QL1 ( .IN(Q0), .IP(P), .IZ(Q2) );

endmodule // ckdpad

`endif

`ifdef bpad8
`else
`define bpad8
module bpad8( A , EN, Q, P );
 input [7:0] A;
input EN;
 inout [7:0] P;
 output [7:0] Q;

bipad QL1 ( .A(A[0]), .EN(EN), .P(P[0]), .Q(Q[0]) );
bipad QL2 ( .A(A[1]), .EN(EN), .P(P[1]), .Q(Q[1]) );
bipad QL3 ( .A(A[2]), .EN(EN), .P(P[2]), .Q(Q[2]) );
bipad QL4 ( .A(A[3]), .EN(EN), .P(P[3]), .Q(Q[3]) );
bipad QL5 ( .A(A[4]), .EN(EN), .P(P[4]), .Q(Q[4]) );
bipad QL6 ( .A(A[5]), .EN(EN), .P(P[5]), .Q(Q[5]) );
bipad QL7 ( .A(A[6]), .EN(EN), .P(P[6]), .Q(Q[6]) );
bipad QL8 ( .A(A[7]), .EN(EN), .P(P[7]), .Q(Q[7]) );

endmodule // bpad8

`endif

`ifdef bpad4
`else
`define bpad4
module bpad4( A , EN, Q, P );
 input [3:0] A;
input EN;
 inout [3:0] P;
 output [3:0] Q;

bipad QL1 ( .A(A[0]), .EN(EN), .P(P[0]), .Q(Q[0]) );
bipad QL2 ( .A(A[1]), .EN(EN), .P(P[1]), .Q(Q[1]) );
bipad QL3 ( .A(A[2]), .EN(EN), .P(P[2]), .Q(Q[2]) );
bipad QL4 ( .A(A[3]), .EN(EN), .P(P[3]), .Q(Q[3]) );

endmodule // bpad4

`endif

`ifdef bpad16
`else
`define bpad16
module bpad16( A , EN, Q, P );
 input [15:0] A;
input EN;
 inout [15:0] P;
 output [15:0] Q;

bipad QL1 ( .A(A[15]), .EN(EN), .P(P[15]), .Q(Q[15]) );
bipad QL2 ( .A(A[14]), .EN(EN), .P(P[14]), .Q(Q[14]) );
bipad QL3 ( .A(A[13]), .EN(EN), .P(P[13]), .Q(Q[13]) );
bipad QL4 ( .A(A[12]), .EN(EN), .P(P[12]), .Q(Q[12]) );
bipad QL5 ( .A(A[11]), .EN(EN), .P(P[11]), .Q(Q[11]) );
bipad QL6 ( .A(A[10]), .EN(EN), .P(P[10]), .Q(Q[10]) );
bipad QL7 ( .A(A[9]), .EN(EN), .P(P[9]), .Q(Q[9]) );
bipad QL8 ( .A(A[8]), .EN(EN), .P(P[8]), .Q(Q[8]) );
bipad QL9 ( .A(A[7]), .EN(EN), .P(P[7]), .Q(Q[7]) );
bipad QL10 ( .A(A[6]), .EN(EN), .P(P[6]), .Q(Q[6]) );
bipad QL11 ( .A(A[5]), .EN(EN), .P(P[5]), .Q(Q[5]) );
bipad QL12 ( .A(A[4]), .EN(EN), .P(P[4]), .Q(Q[4]) );
bipad QL13 ( .A(A[3]), .EN(EN), .P(P[3]), .Q(Q[3]) );
bipad QL14 ( .A(A[2]), .EN(EN), .P(P[2]), .Q(Q[2]) );
bipad QL15 ( .A(A[1]), .EN(EN), .P(P[1]), .Q(Q[1]) );
bipad QL16 ( .A(A[0]), .EN(EN), .P(P[0]), .Q(Q[0]) );

endmodule // bpad16

`endif

`ifdef bipados
`else
`define bipados
module bipados( EN , Q, P );
input EN;
inout P;
output Q;
parameter ql_gate = `BIDIR;
supply1 VCC;
supply0 GND;

bicell QL1 ( .I1(GND), .I2(VCC), .IE(EN), .IP(P), .IZ(Q) );

endmodule // bipados

`endif

`ifdef bipadod
`else
`define bipadod
module bipadod( EN , Q, P );
input EN;
inout P;
output Q;
parameter ql_gate = `BIDIR;
supply1 VCC;
supply0 GND;

bicell QL1 ( .I1(VCC), .I2(GND), .IE(EN), .IP(P), .IZ(Q) );

endmodule // bipadod

`endif

`ifdef bipad
`else
`define bipad
module bipad( A , EN, Q, P );
input A, EN;
inout P;
output Q;
parameter ql_gate = `BIDIR;
supply1 VCC;

bicell QL1 ( .I1(VCC), .I2(A), .IE(EN), .IP(P), .IZ(Q) );

endmodule // bipad

`endif

`ifdef biorpad
`else
`define biorpad
module biorpad( A1 , A2, EN, Q, P );
input A1, A2, EN;
inout P;
output Q;
parameter ql_gate = `BIDIR;

bicell QL1 ( .I1(A1), .I2(A2), .IE(EN), .IP(P), .IZ(Q) );

endmodule // biorpad

`endif

`ifdef biipad
`else
`define biipad
module biipad( A , EN, Q, P );
input A, EN;
inout P;
output Q;
parameter ql_gate = `BIDIR;
supply0 GND;

bicell QL1 ( .I1(A), .I2(GND), .IE(EN), .IP(P), .IZ(Q) );

endmodule // biipad

`endif

`ifdef xor3i0
`else
`define xor3i0
module xor3i0( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
supply0 GND;
supply1 VCC;
wire N_1;
wire N_2;

frag_m I_2 ( .B1(C), .B2(GND), .C1(VCC), .C2(C), .D1(VCC), .D2(C), .E1(C), .E2(GND),
          .NS(N_2), .OS(N_1), .OZ(Q) );
frag_f I_1 ( .F1(B), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );
frag_a QL1 ( .A1(A), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_1) );

endmodule // xor3i0

`endif

`ifdef xor2i0
`else
`define xor2i0
module xor2i0( A , B, Q );
input A, B;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
supply1 VCC;
wire N_2;

frag_a I_2 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(B), .D2(GND), .E1(VCC),
          .E2(B), .NS(N_2), .NZ(Q), .OS(N_1) );
frag_f QL1 ( .F1(A), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );

endmodule // xor2i0

`endif

`ifdef xnor3i0
`else
`define xnor3i0
module xnor3i0( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
supply0 GND;
supply1 VCC;
wire N_1;
wire N_2;

frag_m I_2 ( .B1(VCC), .B2(C), .C1(C), .C2(GND), .D1(C), .D2(GND), .E1(VCC), .E2(C),
          .NS(N_2), .OS(N_1), .OZ(Q) );
frag_f I_1 ( .F1(B), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );
frag_a QL1 ( .A1(A), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_1) );

endmodule // xnor3i0

`endif

`ifdef xnor2i0
`else
`define xnor2i0
module xnor2i0( A , B, Q );
input A, B;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
supply1 VCC;
wire N_2;

frag_a I_2 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(B), .E1(B),
          .E2(GND), .NS(N_2), .NZ(Q), .OS(N_1) );
frag_f QL1 ( .F1(A), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );

endmodule // xnor2i0

`endif

`ifdef sop14i7
`else
`define sop14i7
module sop14i7( A , B, C, D, E, F, G, H, I, J, K, L, M, N, Q );
input A, B, C, D, E, F, G, H, I, J, K, L, M, N;
output Q;
parameter ql_gate = `LOGIC;
supply0 GND;
supply1 VCC;
wire N_1;
wire N_2;

frag_m I_2 ( .B1(G), .B2(H), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(VCC),
          .E2(GND), .NS(N_2), .OS(N_1), .OZ(Q) );
frag_f I_1 ( .F1(I), .F2(L), .F3(J), .F4(M), .F5(K), .F6(N), .FZ(N_2) );
frag_a QL1 ( .A1(A), .A2(D), .A3(B), .A4(E), .A5(C), .A6(F), .AZ(N_1) );

endmodule // sop14i7

`endif

`ifdef maj3i0
`else
`define maj3i0
module maj3i0( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
supply0 GND;
supply1 VCC;
wire N_1;
wire N_2;

frag_m I_2 ( .B1(GND), .B2(VCC), .C1(C), .C2(GND), .D1(C), .D2(GND), .E1(VCC),
          .E2(GND), .NS(N_2), .OS(N_1), .OZ(Q) );
frag_f I_1 ( .F1(B), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );
frag_a QL1 ( .A1(A), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_1) );

endmodule // maj3i0

`endif

`ifdef logicq
`else
`define logicq
module logicq( QC , QD, QR, QS, QZ );
input QC, QR, QS, QD;
output QZ;

p_ff QL1 ( .C(QC), .D(QD), .Q(QZ), .R(QR), .S(QS) );

endmodule // logicq

`endif

`ifdef logicm
`else
`define logicm
module logicm( B1 , B2, C1, C2, D1, D2, E1, E2, NS, OS, NZ, OZ );
input B1, B2, C1, C2, D1, D2, E1, E2, NS;
output NZ;
input OS;
output OZ;

p_mux3 QL2 ( .A(B1), .B(B2), .C(C1), .D(C2), .E(NZ), .S(NS), .T(OS), .Z(OZ) );
p_mux2 QL1 ( .A(D1), .B(D2), .C(E1), .D(E2), .S(NS), .Z(NZ) );

endmodule // logicm

`endif

`ifdef logicf
`else
`define logicf
module logicf( F1 , F2, F3, F4, F5, F6, FZ );
input F1, F2, F3, F4, F5, F6;
output FZ;

p_and6 QL1 ( .A(F1), .B(F2), .C(F3), .D(F4), .E(F5), .F(F6), .Z(FZ) );

endmodule // logicf

`endif

`ifdef logica
`else
`define logica
module logica( A1 , A2, A3, A4, A5, A6, AZ );
input A1, A2, A3, A4, A5, A6;
output AZ;

p_and6 QL1 ( .A(A1), .B(A2), .C(A3), .D(A4), .E(A5), .F(A6), .Z(AZ) );

endmodule // logica

`endif

`ifdef inv
`else
`define inv
module inv( A , Q );
input A;
output Q;
supply1 VCC;

nand2i0 I1 ( .A(VCC), .B(A), .Q(Q) );

endmodule // inv

`endif

`ifdef dece2t4
`else
`define dece2t4
module dece2t4( EN , S0, S1, Q0, Q1, Q2, Q3 );
input EN;
output Q0, Q1, Q2, Q3;
input S0, S1;

and3i0 QL1 ( .A(EN), .B(S0), .C(S1), .Q(Q3) );
and3i1 QL2 ( .A(EN), .B(S1), .C(S0), .Q(Q2) );
and3i1 QL3 ( .A(EN), .B(S0), .C(S1), .Q(Q1) );
and3i2 QL4 ( .A(EN), .B(S0), .C(S1), .Q(Q0) );

endmodule // dece2t4

`endif

`ifdef dec2t4
`else
`define dec2t4
module dec2t4( S0 , S1, Q0, Q1, Q2, Q3 );
output Q0, Q1, Q2, Q3;
input S0, S1;
parameter ql_gate = `LOGIC;
supply0 GND;
supply1 VCC;

frag_m I_2 ( .B1(S0), .B2(S1), .C1(GND), .C2(VCC), .D1(S1), .D2(S0), .E1(GND),
          .E2(VCC), .NS(Q3), .NZ(Q2), .OS(Q0), .OZ(Q1) );
frag_f I_1 ( .F1(S0), .F2(GND), .F3(S1), .F4(GND), .F5(VCC), .F6(GND), .FZ(Q3) );
frag_a QL1 ( .A1(VCC), .A2(S0), .A3(VCC), .A4(S1), .A5(VCC), .A6(GND), .AZ(Q0) );

endmodule // dec2t4

`endif

`ifdef buff
`else
`define buff
module buff( A , Q );
input A;
output Q;
parameter ql_gate = `LOGIC;
supply0 GND;
supply1 VCC;

frag_a QL1 ( .A1(A), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(Q) );

endmodule // buff

`endif

`ifdef or6i6
`else
`define or6i6
module or6i6( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(D), .A2(GND), .A3(E), .A4(GND), .A5(F), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(A), .F2(GND), .F3(B), .F4(GND), .F5(C), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // or6i6

`endif

`ifdef or6i5
`else
`define or6i5
module or6i5( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(D), .A2(GND), .A3(E), .A4(GND), .A5(F), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(VCC), .F2(A), .F3(B), .F4(GND), .F5(C), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // or6i5

`endif

`ifdef or6i4
`else
`define or6i4
module or6i4( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(D), .F2(A), .F3(E), .F4(B), .F5(F), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(VCC),
          .E2(C), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or6i4

`endif

`ifdef or6i3
`else
`define or6i3
module or6i3( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(D), .F2(A), .F3(E), .F4(B), .F5(F), .F6(C), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or6i3

`endif

`ifdef or6i2
`else
`define or6i2
module or6i2( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(VCC), .F2(A), .F3(E), .F4(B), .F5(F), .F6(C), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(D),
          .E2(GND), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or6i2

`endif

`ifdef or6i1
`else
`define or6i1
module or6i1( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(VCC), .A2(D), .A3(VCC), .A4(E), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(F), .F6(C), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // or6i1

`endif

`ifdef or6i0
`else
`define or6i0
module or6i0( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(VCC), .A2(D), .A3(VCC), .A4(E), .A5(VCC), .A6(F), .AZ(N_2) );
frag_f I_1 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // or6i0

`endif

`ifdef or5i5
`else
`define or5i5
module or5i5( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(D), .A2(GND), .A3(E), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(A), .F2(GND), .F3(B), .F4(GND), .F5(C), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // or5i5

`endif

`ifdef or5i4
`else
`define or5i4
module or5i4( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(C), .F2(A), .F3(D), .F4(GND), .F5(E), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(VCC),
          .E2(B), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or5i4

`endif

`ifdef or5i3
`else
`define or5i3
module or5i3( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(D), .F2(A), .F3(E), .F4(B), .F5(C), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or5i3

`endif

`ifdef or5i2
`else
`define or5i2
module or5i2( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(VCC), .F2(A), .F3(D), .F4(B), .F5(E), .F6(C), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or5i2

`endif

`ifdef or5i1
`else
`define or5i1
module or5i1( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(E), .F6(C), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(D),
          .E2(GND), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or5i1

`endif

`ifdef or5i0
`else
`define or5i0
module or5i0( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(VCC), .A2(D), .A3(VCC), .A4(E), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // or5i0

`endif

`ifdef or4i4
`else
`define or4i4
module or4i4( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(B), .F2(GND), .F3(C), .F4(GND), .F5(D), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(VCC),
          .E2(A), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or4i4

`endif

`ifdef or4i3
`else
`define or4i3
module or4i3( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(D), .F2(A), .F3(B), .F4(GND), .F5(C), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or4i3

`endif

`ifdef or4i2
`else
`define or4i2
module or4i2( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(VCC), .F2(A), .F3(D), .F4(B), .F5(C), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or4i2

`endif

`ifdef or4i1
`else
`define or4i1
module or4i1( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(VCC), .F2(A), .F3(D), .F4(B), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or4i1

`endif

`ifdef or4i0
`else
`define or4i0
module or4i0( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(D),
          .E2(GND), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or4i0

`endif

`ifdef or3i3
`else
`define or3i3
module or3i3( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(A), .F2(GND), .F3(B), .F4(GND), .F5(C), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or3i3

`endif

`ifdef or3i2
`else
`define or3i2
module or3i2( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(VCC), .F2(A), .F3(B), .F4(GND), .F5(C), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or3i2

`endif

`ifdef or3i1
`else
`define or3i1
module or3i1( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(C), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or3i1

`endif

`ifdef or3i0
`else
`define or3i0
module or3i0( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or3i0

`endif

`ifdef or2i2
`else
`define or2i2
module or2i2( A , B, Q );
input A, B;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(A), .F2(GND), .F3(B), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or2i2

`endif

`ifdef or2i1
`else
`define or2i1
module or2i1( A , B, Q );
input A, B;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(VCC), .F2(A), .F3(B), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or2i1

`endif

`ifdef or2i0
`else
`define or2i0
module or2i0( A , B, Q );
input A, B;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // or2i0

`endif

`ifdef or13i6
`else
`define or13i6
module or13i6( A , B, C, D, E, F, G, H, I, J, K, L, M, Q );
input A, B, C, D, E, F, G, H, I, J, K, L, M;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(H), .A2(A), .A3(I), .A4(B), .A5(J), .A6(C), .AZ(N_2) );
frag_f I_1 ( .F1(K), .F2(E), .F3(L), .F4(F), .F5(M), .F6(G), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(D),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // or13i6

`endif

`ifdef nor6i6
`else
`define nor6i6
module nor6i6( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(D), .A2(GND), .A3(E), .A4(GND), .A5(F), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(A), .F2(GND), .F3(B), .F4(GND), .F5(C), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(GND), .B2(VCC), .C1(GND), .C2(VCC), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // nor6i6

`endif

`ifdef nor6i5
`else
`define nor6i5
module nor6i5( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(D), .A2(GND), .A3(E), .A4(GND), .A5(F), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(VCC), .F2(A), .F3(B), .F4(GND), .F5(C), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(GND), .B2(VCC), .C1(GND), .C2(VCC), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // nor6i5

`endif

`ifdef nor6i4
`else
`define nor6i4
module nor6i4( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(D), .F2(A), .F3(E), .F4(B), .F5(F), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(GND), .D2(VCC), .E1(C),
          .E2(GND), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nor6i4

`endif

`ifdef nor6i3
`else
`define nor6i3
module nor6i3( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;

frag_a QL1 ( .A1(D), .A2(A), .A3(E), .A4(B), .A5(F), .A6(C), .AZ(Q) );

endmodule // nor6i3

`endif

`ifdef nor6i2
`else
`define nor6i2
module nor6i2( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(VCC), .F2(A), .F3(E), .F4(B), .F5(F), .F6(C), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(D), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nor6i2

`endif

`ifdef nor6i1
`else
`define nor6i1
module nor6i1( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(VCC), .A2(D), .A3(VCC), .A4(E), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(F), .F6(C), .FZ(N_1) );
frag_m QL3 ( .B1(GND), .B2(VCC), .C1(GND), .C2(VCC), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // nor6i1

`endif

`ifdef nor6i0
`else
`define nor6i0
module nor6i0( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(VCC), .A2(D), .A3(VCC), .A4(E), .A5(VCC), .A6(F), .AZ(N_2) );
frag_f I_1 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m QL3 ( .B1(GND), .B2(VCC), .C1(GND), .C2(VCC), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // nor6i0

`endif

`ifdef nor5i5
`else
`define nor5i5
module nor5i5( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(D), .A2(GND), .A3(E), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(A), .F2(GND), .F3(B), .F4(GND), .F5(C), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(GND), .B2(VCC), .C1(GND), .C2(VCC), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // nor5i5

`endif

`ifdef nor5i4
`else
`define nor5i4
module nor5i4( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(C), .F2(A), .F3(D), .F4(GND), .F5(E), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(GND), .D2(VCC), .E1(B),
          .E2(GND), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nor5i4

`endif

`ifdef nor5i3
`else
`define nor5i3
module nor5i3( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
supply0 GND;

frag_a QL1 ( .A1(D), .A2(GND), .A3(E), .A4(A), .A5(C), .A6(B), .AZ(Q) );

endmodule // nor5i3

`endif

`ifdef nor5i2
`else
`define nor5i2
module nor5i2( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;

frag_a QL1 ( .A1(D), .A2(A), .A3(E), .A4(B), .A5(VCC), .A6(C), .AZ(Q) );

endmodule // nor5i2

`endif

`ifdef nor5i1
`else
`define nor5i1
module nor5i1( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(E), .F6(C), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(D), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nor5i1

`endif

`ifdef nor5i0
`else
`define nor5i0
module nor5i0( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(VCC), .A2(D), .A3(VCC), .A4(E), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m QL3 ( .B1(GND), .B2(VCC), .C1(GND), .C2(VCC), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // nor5i0

`endif

`ifdef nor4i4
`else
`define nor4i4
module nor4i4( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(B), .F2(GND), .F3(C), .F4(GND), .F5(D), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(GND), .D2(VCC), .E1(A),
          .E2(GND), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nor4i4

`endif

`ifdef nor4i3
`else
`define nor4i3
module nor4i3( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
supply0 GND;

frag_a QL1 ( .A1(D), .A2(GND), .A3(B), .A4(GND), .A5(C), .A6(A), .AZ(Q) );

endmodule // nor4i3

`endif

`ifdef nor4i2
`else
`define nor4i2
module nor4i2( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

frag_a QL1 ( .A1(D), .A2(GND), .A3(C), .A4(A), .A5(VCC), .A6(B), .AZ(Q) );

endmodule // nor4i2

`endif

`ifdef nor4i1
`else
`define nor4i1
module nor4i1( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;

frag_a QL1 ( .A1(D), .A2(A), .A3(VCC), .A4(B), .A5(VCC), .A6(C), .AZ(Q) );

endmodule // nor4i1

`endif

`ifdef nor4i0
`else
`define nor4i0
module nor4i0( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(D), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nor4i0

`endif

`ifdef nor3i3
`else
`define nor3i3
module nor3i3( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
supply0 GND;

frag_a QL1 ( .A1(A), .A2(GND), .A3(B), .A4(GND), .A5(C), .A6(GND), .AZ(Q) );

endmodule // nor3i3

`endif

`ifdef nor3i2
`else
`define nor3i2
module nor3i2( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

frag_a QL1 ( .A1(B), .A2(GND), .A3(C), .A4(GND), .A5(VCC), .A6(A), .AZ(Q) );

endmodule // nor3i2

`endif

`ifdef nor3i1
`else
`define nor3i1
module nor3i1( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

frag_a QL1 ( .A1(C), .A2(GND), .A3(VCC), .A4(A), .A5(VCC), .A6(B), .AZ(Q) );

endmodule // nor3i1

`endif

`ifdef nor3i0
`else
`define nor3i0
module nor3i0( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;

frag_a QL1 ( .A1(VCC), .A2(A), .A3(VCC), .A4(B), .A5(VCC), .A6(C), .AZ(Q) );

endmodule // nor3i0

`endif

`ifdef nor2i2
`else
`define nor2i2
module nor2i2( A , B, Q );
input A, B;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

frag_a QL1 ( .A1(A), .A2(GND), .A3(B), .A4(GND), .A5(VCC), .A6(GND), .AZ(Q) );

endmodule // nor2i2

`endif

`ifdef nor2i1
`else
`define nor2i1
module nor2i1( A , B, Q );
input A, B;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

frag_a QL1 ( .A1(B), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(A), .AZ(Q) );

endmodule // nor2i1

`endif

`ifdef nor2i0
`else
`define nor2i0
module nor2i0( A , B, Q );
input A, B;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

frag_a QL1 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(A), .A5(VCC), .A6(B), .AZ(Q) );

endmodule // nor2i0

`endif

`ifdef nor14i7
`else
`define nor14i7
module nor14i7( A , B, C, D, E, F, G, H, I, J, K, L, M, N, Q );
input A, B, C, D, E, F, G, H, I, J, K, L, M, N;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(H), .A2(A), .A3(I), .A4(B), .A5(J), .A6(C), .AZ(N_2) );
frag_f I_1 ( .F1(L), .F2(E), .F3(M), .F4(F), .F5(N), .F6(G), .FZ(N_1) );
frag_m QL3 ( .B1(GND), .B2(VCC), .C1(GND), .C2(VCC), .D1(GND), .D2(VCC), .E1(K),
          .E2(D), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // nor14i7

`endif

`ifdef nand6i6
`else
`define nand6i6
module nand6i6( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(VCC), .A2(D), .A3(VCC), .A4(E), .A5(VCC), .A6(F), .AZ(N_2) );
frag_f I_1 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // nand6i6

`endif

`ifdef nand6i5
`else
`define nand6i5
module nand6i5( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(VCC), .A2(D), .A3(VCC), .A4(E), .A5(VCC), .A6(F), .AZ(N_2) );
frag_f I_1 ( .F1(A), .F2(GND), .F3(VCC), .F4(B), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // nand6i5

`endif

`ifdef nand6i4
`else
`define nand6i4
module nand6i4( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(A), .F2(D), .F3(B), .F4(E), .F5(VCC), .F6(F), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(C),
          .E2(GND), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand6i4

`endif

`ifdef nand6i3
`else
`define nand6i3
module nand6i3( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(A), .F2(D), .F3(B), .F4(E), .F5(C), .F6(F), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand6i3

`endif

`ifdef nand6i2
`else
`define nand6i2
module nand6i2( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(A), .F2(GND), .F3(B), .F4(E), .F5(C), .F6(F), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(VCC),
          .E2(D), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand6i2

`endif

`ifdef nand6i1
`else
`define nand6i1
module nand6i1( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(D), .A2(GND), .A3(E), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(A), .F2(GND), .F3(B), .F4(GND), .F5(C), .F6(F), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // nand6i1

`endif

`ifdef nand6i0
`else
`define nand6i0
module nand6i0( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(D), .A2(GND), .A3(E), .A4(GND), .A5(F), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(A), .F2(GND), .F3(B), .F4(GND), .F5(C), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // nand6i0

`endif

`ifdef nand5i5
`else
`define nand5i5
module nand5i5( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(VCC), .A2(D), .A3(VCC), .A4(E), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // nand5i5

`endif

`ifdef nand5i4
`else
`define nand5i4
module nand5i4( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(A), .F2(C), .F3(VCC), .F4(D), .F5(VCC), .F6(E), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(B),
          .E2(GND), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand5i4

`endif

`ifdef nand5i3
`else
`define nand5i3
module nand5i3( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(A), .F2(D), .F3(B), .F4(E), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand5i3

`endif

`ifdef nand5i2
`else
`define nand5i2
module nand5i2( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(A), .F2(D), .F3(B), .F4(E), .F5(C), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand5i2

`endif

`ifdef nand5i1
`else
`define nand5i1
module nand5i1( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(A), .F2(GND), .F3(B), .F4(E), .F5(C), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(VCC),
          .E2(D), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand5i1

`endif

`ifdef nand5i0
`else
`define nand5i0
module nand5i0( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(D), .A2(GND), .A3(E), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(A), .F2(GND), .F3(B), .F4(GND), .F5(C), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // nand5i0

`endif

`ifdef nand4i4
`else
`define nand4i4
module nand4i4( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(VCC), .F2(B), .F3(VCC), .F4(C), .F5(VCC), .F6(D), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(A),
          .E2(GND), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand4i4

`endif

`ifdef nand4i3
`else
`define nand4i3
module nand4i3( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(A), .F2(D), .F3(VCC), .F4(B), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand4i3

`endif

`ifdef nand4i2
`else
`define nand4i2
module nand4i2( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(A), .F2(D), .F3(B), .F4(GND), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand4i2

`endif

`ifdef nand4i1
`else
`define nand4i1
module nand4i1( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(A), .F2(D), .F3(B), .F4(GND), .F5(C), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand4i1

`endif

`ifdef nand4i0
`else
`define nand4i0
module nand4i0( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(A), .F2(GND), .F3(B), .F4(GND), .F5(C), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(VCC),
          .E2(D), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand4i0

`endif

`ifdef nand3i3
`else
`define nand3i3
module nand3i3( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand3i3

`endif

`ifdef nand3i2
`else
`define nand3i2
module nand3i2( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(A), .F2(GND), .F3(VCC), .F4(B), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand3i2

`endif

`ifdef nand3i1
`else
`define nand3i1
module nand3i1( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(A), .F2(GND), .F3(B), .F4(GND), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand3i1

`endif

`ifdef nand3i0
`else
`define nand3i0
module nand3i0( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(A), .F2(GND), .F3(B), .F4(GND), .F5(C), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand3i0

`endif

`ifdef nand2i2
`else
`define nand2i2
module nand2i2( A , B, Q );
input A, B;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand2i2

`endif

`ifdef nand2i1
`else
`define nand2i1
module nand2i1( A , B, Q );
input A, B;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(A), .F2(GND), .F3(VCC), .F4(B), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand2i1

`endif

`ifdef nand2i0
`else
`define nand2i0
module nand2i0( A , B, Q );
input A, B;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(A), .F2(GND), .F3(B), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // nand2i0

`endif

`ifdef nand13i6
`else
`define nand13i6
module nand13i6( A , B, C, D, E, F, G, H, I, J, K, L, M, Q );
input A, B, C, D, E, F, G, H, I, J, K, L, M;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(A), .A2(H), .A3(B), .A4(I), .A5(C), .A6(J), .AZ(N_2) );
frag_f I_1 ( .F1(E), .F2(K), .F3(F), .F4(L), .F5(G), .F6(M), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(VCC),
          .E2(D), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // nand13i6

`endif

`ifdef mux4xf
`else
`define mux4xf
module mux4xf( A , B, C, D, S0, S1, Q );
input A, B, C, D;
output Q;
input S0, S1;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(A), .C1(VCC), .C2(B), .D1(VCC), .D2(C), .E1(VCC), .E2(D),
          .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // mux4xf

`endif

`ifdef mux4xe
`else
`define mux4xe
module mux4xe( A , B, C, D, S0, S1, Q );
input A, B, C, D;
output Q;
input S0, S1;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(A), .B2(GND), .C1(VCC), .C2(B), .D1(VCC), .D2(C), .E1(VCC), .E2(D),
          .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // mux4xe

`endif

`ifdef mux4xd
`else
`define mux4xd
module mux4xd( A , B, C, D, S0, S1, Q );
input A, B, C, D;
output Q;
input S0, S1;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(A), .C1(B), .C2(GND), .D1(VCC), .D2(C), .E1(VCC), .E2(D),
          .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // mux4xd

`endif

`ifdef mux4xc
`else
`define mux4xc
module mux4xc( A , B, C, D, S0, S1, Q );
input A, B, C, D;
output Q;
input S0, S1;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(A), .B2(GND), .C1(B), .C2(GND), .D1(VCC), .D2(C), .E1(VCC), .E2(D),
          .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // mux4xc

`endif

`ifdef mux4xb
`else
`define mux4xb
module mux4xb( A , B, C, D, S0, S1, Q );
input A, B, C, D;
output Q;
input S0, S1;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(A), .C1(VCC), .C2(B), .D1(C), .D2(GND), .E1(VCC), .E2(D),
          .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // mux4xb

`endif

`ifdef mux4xa
`else
`define mux4xa
module mux4xa( A , B, C, D, S0, S1, Q );
input A, B, C, D;
output Q;
input S0, S1;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(A), .B2(GND), .C1(VCC), .C2(B), .D1(C), .D2(GND), .E1(VCC), .E2(D),
          .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // mux4xa

`endif

`ifdef mux4x9
`else
`define mux4x9
module mux4x9( A , B, C, D, S0, S1, Q );
input A, B, C, D;
output Q;
input S0, S1;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(A), .C1(B), .C2(GND), .D1(C), .D2(GND), .E1(VCC), .E2(D),
          .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // mux4x9

`endif

`ifdef mux4x8
`else
`define mux4x8
module mux4x8( A , B, C, D, S0, S1, Q );
input A, B, C, D;
output Q;
input S0, S1;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(A), .B2(GND), .C1(B), .C2(GND), .D1(C), .D2(GND), .E1(VCC), .E2(D),
          .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // mux4x8

`endif

`ifdef mux4x7
`else
`define mux4x7
module mux4x7( A , B, C, D, S0, S1, Q );
input A, B, C, D;
output Q;
input S0, S1;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(A), .C1(VCC), .C2(B), .D1(VCC), .D2(C), .E1(D), .E2(GND),
          .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // mux4x7

`endif

`ifdef mux4x6
`else
`define mux4x6
module mux4x6( A , B, C, D, S0, S1, Q );
input A, B, C, D;
output Q;
input S0, S1;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(A), .B2(GND), .C1(VCC), .C2(B), .D1(VCC), .D2(C), .E1(D), .E2(GND),
          .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // mux4x6

`endif

`ifdef mux4x5
`else
`define mux4x5
module mux4x5( A , B, C, D, S0, S1, Q );
input A, B, C, D;
output Q;
input S0, S1;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(A), .C1(B), .C2(GND), .D1(VCC), .D2(C), .E1(D), .E2(GND),
          .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // mux4x5

`endif

`ifdef mux4x4
`else
`define mux4x4
module mux4x4( A , B, C, D, S0, S1, Q );
input A, B, C, D;
output Q;
input S0, S1;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(A), .B2(GND), .C1(B), .C2(GND), .D1(VCC), .D2(C), .E1(D), .E2(GND),
          .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // mux4x4

`endif

`ifdef mux4x3
`else
`define mux4x3
module mux4x3( A , B, C, D, S0, S1, Q );
input A, B, C, D;
output Q;
input S0, S1;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(A), .C1(VCC), .C2(B), .D1(C), .D2(GND), .E1(D), .E2(GND),
          .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // mux4x3

`endif

`ifdef mux4x2
`else
`define mux4x2
module mux4x2( A , B, C, D, S0, S1, Q );
input A, B, C, D;
output Q;
input S0, S1;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(A), .B2(GND), .C1(VCC), .C2(B), .D1(C), .D2(GND), .E1(D), .E2(GND),
          .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // mux4x2

`endif

`ifdef mux4x1
`else
`define mux4x1
module mux4x1( A , B, C, D, S0, S1, Q );
input A, B, C, D;
output Q;
input S0, S1;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(VCC), .B2(A), .C1(B), .C2(GND), .D1(C), .D2(GND), .E1(D), .E2(GND),
          .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // mux4x1

`endif

`ifdef mux4x0
`else
`define mux4x0
module mux4x0( A , B, C, D, S0, S1, Q );
input A, B, C, D;
output Q;
input S0, S1;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(A), .B2(GND), .C1(B), .C2(GND), .D1(C), .D2(GND), .E1(D), .E2(GND),
          .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // mux4x0

`endif

`ifdef mux2x3
`else
`define mux2x3
module mux2x3( A , B, S, Q );
input A, B;
output Q;
input S;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(S), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(A), .E1(VCC),
          .E2(B), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // mux2x3

`endif

`ifdef mux2x2
`else
`define mux2x2
module mux2x2( A , B, S, Q );
input A, B;
output Q;
input S;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(S), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(A), .D2(GND), .E1(VCC),
          .E2(B), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // mux2x2

`endif

`ifdef mux2x1
`else
`define mux2x1
module mux2x1( A , B, S, Q );
input A, B;
output Q;
input S;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(S), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(A), .E1(B),
          .E2(GND), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // mux2x1

`endif

`ifdef mux2x0
`else
`define mux2x0
module mux2x0( A , B, S, Q );
input A, B;
output Q;
input S;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(S), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(A), .D2(GND), .E1(B),
          .E2(GND), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // mux2x0

`endif

`ifdef mux2ffx3
`else
`define mux2ffx3
module mux2ffx3( A , CLK, CLR, D, PRE, S, Q, R );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input PRE /* synthesis syn_isclock=1 */;
input A, D;
output Q, R;
input S;
parameter syn_macro = 1, ql_pack = 1;
parameter ql_gate = `LOGIC;
supply0 GND;
wire N_1;
supply1 VCC;
wire N_2;
wire N_3;

frag_m I_3 ( .B1(D), .B2(GND), .C1(D), .C2(GND), .D1(VCC), .D2(A), .E1(VCC), .E2(Q),
          .NS(N_3), .NZ(R), .OS(N_2), .OZ(N_1) );
frag_q I_2 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(PRE), .QZ(Q) );
frag_a I_1 ( .A1(GND), .A2(VCC), .A3(GND), .A4(VCC), .A5(GND), .A6(VCC), .AZ(N_2) );
frag_f QL4 ( .F1(S), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_3) );

endmodule // mux2ffx3

`endif

`ifdef mux2ffx2
`else
`define mux2ffx2
module mux2ffx2( A , CLK, CLR, D, PRE, S, Q, R );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input PRE /* synthesis syn_isclock=1 */;
input A, D;
output Q, R;
input S;
parameter syn_macro = 1, ql_pack = 1;
parameter ql_gate = `LOGIC;
supply0 GND;
wire N_1;
supply1 VCC;
wire N_2;
wire N_3;

frag_m I_3 ( .B1(D), .B2(GND), .C1(D), .C2(GND), .D1(A), .D2(GND), .E1(VCC), .E2(Q),
          .NS(N_3), .NZ(R), .OS(N_2), .OZ(N_1) );
frag_q I_2 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(PRE), .QZ(Q) );
frag_a I_1 ( .A1(GND), .A2(VCC), .A3(GND), .A4(VCC), .A5(GND), .A6(VCC), .AZ(N_2) );
frag_f QL4 ( .F1(S), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_3) );

endmodule // mux2ffx2

`endif

`ifdef mux2ffx1
`else
`define mux2ffx1
module mux2ffx1( A , CLK, CLR, D, PRE, S, Q, R );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input PRE /* synthesis syn_isclock=1 */;
input A, D;
output Q, R;
input S;
parameter syn_macro = 1, ql_pack = 1;
parameter ql_gate = `LOGIC;
supply0 GND;
wire N_1;
supply1 VCC;
wire N_2;
wire N_3;

frag_m I_3 ( .B1(D), .B2(GND), .C1(D), .C2(GND), .D1(VCC), .D2(A), .E1(Q), .E2(GND),
          .NS(N_3), .NZ(R), .OS(N_2), .OZ(N_1) );
frag_q I_2 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(PRE), .QZ(Q) );
frag_a I_1 ( .A1(GND), .A2(VCC), .A3(GND), .A4(VCC), .A5(GND), .A6(VCC), .AZ(N_2) );
frag_f QL4 ( .F1(S), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_3) );

endmodule // mux2ffx1

`endif

`ifdef mux2ffx0
`else
`define mux2ffx0
module mux2ffx0( A , CLK, CLR, D, PRE, S, Q, R );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input PRE /* synthesis syn_isclock=1 */;
input A, D;
output Q, R;
input S;
parameter syn_macro = 1, ql_pack = 1;
parameter ql_gate = `LOGIC;
supply0 GND;
wire N_1;
supply1 VCC;
wire N_2;
wire N_3;

frag_m I_3 ( .B1(D), .B2(GND), .C1(D), .C2(GND), .D1(A), .D2(GND), .E1(Q), .E2(GND),
          .NS(N_3), .NZ(R), .OS(N_2), .OZ(N_1) );
frag_q I_2 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(PRE), .QZ(Q) );
frag_a I_1 ( .A1(GND), .A2(VCC), .A3(GND), .A4(VCC), .A5(GND), .A6(VCC), .AZ(N_2) );
frag_f QL4 ( .F1(S), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_3) );

endmodule // mux2ffx0

`endif

`ifdef mux2dx3
`else
`define mux2dx3
module mux2dx3( A , B, C, D, S, Q, R );
input A, B, C, D;
output Q, R;
input S;
parameter syn_macro = 1, ql_pack = 1;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;
wire N_1;
wire N_2;

frag_a I_2 ( .A1(GND), .A2(VCC), .A3(GND), .A4(VCC), .A5(GND), .A6(VCC), .AZ(N_1) );
frag_f I_1 ( .F1(S), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );
frag_m QL3 ( .B1(VCC), .B2(A), .C1(VCC), .C2(B), .D1(VCC), .D2(C), .E1(VCC), .E2(D),
          .NS(N_2), .NZ(R), .OS(N_1), .OZ(Q) );

endmodule // mux2dx3

`endif

`ifdef mux2dx2
`else
`define mux2dx2
module mux2dx2( A , B, C, D, S, Q, R );
input A, B, C, D;
output Q, R;
input S;
parameter syn_macro = 1, ql_pack = 1;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;
wire N_1;
wire N_2;

frag_a I_2 ( .A1(GND), .A2(VCC), .A3(GND), .A4(VCC), .A5(GND), .A6(VCC), .AZ(N_1) );
frag_f I_1 ( .F1(S), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );
frag_m QL3 ( .B1(A), .B2(GND), .C1(VCC), .C2(B), .D1(C), .D2(GND), .E1(VCC), .E2(D),
          .NS(N_2), .NZ(R), .OS(N_1), .OZ(Q) );

endmodule // mux2dx2

`endif

`ifdef mux2dx1
`else
`define mux2dx1
module mux2dx1( A , B, C, D, S, Q, R );
input A, B, C, D;
output Q, R;
input S;
parameter syn_macro = 1, ql_pack = 1;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;
wire N_1;
wire N_2;

frag_a I_2 ( .A1(GND), .A2(VCC), .A3(GND), .A4(VCC), .A5(GND), .A6(VCC), .AZ(N_1) );
frag_f I_1 ( .F1(S), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );
frag_m QL3 ( .B1(VCC), .B2(A), .C1(B), .C2(GND), .D1(VCC), .D2(C), .E1(D), .E2(GND),
          .NS(N_2), .NZ(R), .OS(N_1), .OZ(Q) );

endmodule // mux2dx1

`endif

`ifdef mux2dx0
`else
`define mux2dx0
module mux2dx0( A , B, C, D, S, Q, R );
input A, B, C, D;
output Q, R;
input S;
parameter syn_macro = 1, ql_pack = 1;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;
wire N_1;
wire N_2;

frag_a I_2 ( .A1(GND), .A2(VCC), .A3(GND), .A4(VCC), .A5(GND), .A6(VCC), .AZ(N_1) );
frag_f I_1 ( .F1(S), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );
frag_m QL3 ( .B1(A), .B2(GND), .C1(B), .C2(GND), .D1(C), .D2(GND), .E1(D), .E2(GND),
          .NS(N_2), .NZ(R), .OS(N_1), .OZ(Q) );

endmodule // mux2dx0

`endif

`ifdef dlap
`else
`define dlap
module dlap( D , G, PRE, Q );
input D, G, PRE;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(PRE), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(G), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(Q), .B2(GND), .C1(D), .C2(GND), .D1(VCC), .D2(GND), .E1(VCC),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // dlap

`endif

`ifdef dlamux
`else
`define dlamux
module dlamux( D0 , D1, G, SEL, Q );
input D0, D1, G;
output Q;
input SEL;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(SEL), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(G), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(Q), .B2(GND), .C1(D0), .C2(GND), .D1(Q), .D2(GND), .E1(D1),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // dlamux

`endif

`ifdef dlaemux
`else
`define dlaemux
module dlaemux( D0 , D1, EN, G, SEL, Q );
input D0, D1, EN, G;
output Q;
input SEL;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(SEL), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(G), .F2(GND), .F3(EN), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(Q), .B2(GND), .C1(D0), .C2(GND), .D1(Q), .D2(GND), .E1(D1),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // dlaemux

`endif

`ifdef dlaec
`else
`define dlaec
module dlaec( CLR , D, EN, G, Q );
input CLR, D, EN, G;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(CLR), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(G), .F2(GND), .F3(EN), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(Q), .B2(GND), .C1(D), .C2(GND), .D1(GND), .D2(VCC), .E1(GND),
          .E2(VCC), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // dlaec

`endif

`ifdef dlae
`else
`define dlae
module dlae( D , EN, G, Q );
input D, EN, G;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(G), .F2(GND), .F3(EN), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(Q), .D2(GND), .E1(D),
          .E2(GND), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // dlae

`endif

`ifdef dlade
`else
`define dlade
module dlade( D1 , D2, EN, G, Q1, Q2 );
input D1, D2, EN, G;
output Q1, Q2;
parameter syn_macro = 1, ql_pack = 1;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;
wire N_1;
wire N_2;

frag_a I_2 ( .A1(GND), .A2(VCC), .A3(GND), .A4(VCC), .A5(GND), .A6(VCC), .AZ(N_2) );
frag_f I_1 ( .F1(G), .F2(GND), .F3(EN), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(Q1), .B2(GND), .C1(D1), .C2(GND), .D1(Q2), .D2(GND), .E1(D2),
          .E2(GND), .NS(N_1), .NZ(Q2), .OS(N_2), .OZ(Q1) );

endmodule // dlade

`endif

`ifdef dlad
`else
`define dlad
module dlad( D1 , D2, G, Q1, Q2 );
input D1, D2, G;
output Q1, Q2;
parameter syn_macro = 1, ql_pack = 1;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;
wire N_1;
wire N_2;

frag_a I_2 ( .A1(GND), .A2(VCC), .A3(GND), .A4(VCC), .A5(GND), .A6(VCC), .AZ(N_2) );
frag_f I_1 ( .F1(G), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(Q1), .B2(GND), .C1(D1), .C2(GND), .D1(Q2), .D2(GND), .E1(D2),
          .E2(GND), .NS(N_1), .NZ(Q2), .OS(N_2), .OZ(Q1) );

endmodule // dlad

`endif

`ifdef dlac
`else
`define dlac
module dlac( CLR , D, G, Q );
input CLR, D, G;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(CLR), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(G), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(Q), .B2(GND), .C1(D), .C2(GND), .D1(GND), .D2(VCC), .E1(GND),
          .E2(VCC), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // dlac

`endif

`ifdef dla
`else
`define dla
module dla( D , G, Q );
input D, G;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(G), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(Q), .D2(GND), .E1(D),
          .E2(GND), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // dla

`endif

`ifdef tffpc
`else
`define tffpc
module tffpc( CLK , CLR, PRE, T, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input PRE /* synthesis syn_isclock=1 */;
output Q;
input T;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
wire N_3;
supply0 GND;

frag_a I_3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_1) );
frag_q I_2 ( .QC(CLK), .QD(N_3), .QR(CLR), .QS(PRE), .QZ(Q) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(Q), .D2(GND), .E1(VCC),
          .E2(Q), .NS(N_2), .OS(N_1), .OZ(N_3) );
frag_f QL1 ( .F1(T), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );

endmodule // tffpc

`endif

`ifdef tffepc
`else
`define tffepc
module tffepc( CLK , CLR, EN, PRE, T, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input PRE /* synthesis syn_isclock=1 */;
input EN;
output Q;
input T;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(PRE), .QZ(Q) );
frag_m I_2 ( .B1(Q), .B2(GND), .C1(Q), .C2(GND), .D1(Q), .D2(GND), .E1(VCC), .E2(Q),
          .NS(N_3), .OS(N_2), .OZ(N_1) );
frag_f I_1 ( .F1(T), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_3) );
frag_a QL1 ( .A1(EN), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // tffepc

`endif

`ifdef tffe
`else
`define tffe
module tffe( CLK , EN, T, Q );
input CLK /* synthesis syn_isclock=1 */;
input EN;
output Q;
input T;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(CLK), .QD(N_1), .QR(GND), .QS(GND), .QZ(Q) );
frag_m I_2 ( .B1(Q), .B2(GND), .C1(Q), .C2(GND), .D1(Q), .D2(GND), .E1(VCC), .E2(Q),
          .NS(N_3), .OS(N_2), .OZ(N_1) );
frag_f I_1 ( .F1(T), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_3) );
frag_a QL1 ( .A1(EN), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // tffe

`endif

`ifdef tff
`else
`define tff
module tff( CLK , T, Q );
input CLK /* synthesis syn_isclock=1 */;
output Q;
input T;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
wire N_3;
supply0 GND;

frag_a I_3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_1) );
frag_q I_2 ( .QC(CLK), .QD(N_3), .QR(GND), .QS(GND), .QZ(Q) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(Q), .D2(GND), .E1(VCC),
          .E2(Q), .NS(N_2), .OS(N_1), .OZ(N_3) );
frag_f QL1 ( .F1(T), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );

endmodule // tff

`endif

`ifdef jkffpc
`else
`define jkffpc
module jkffpc( CLK , CLR, J, K, PRE, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input PRE /* synthesis syn_isclock=1 */;
input J, K;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(PRE), .QZ(Q) );
frag_m I_2 ( .B1(Q), .B2(GND), .C1(GND), .C2(VCC), .D1(VCC), .D2(GND), .E1(VCC),
          .E2(Q), .NS(N_3), .OS(N_2), .OZ(N_1) );
frag_f I_1 ( .F1(K), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_3) );
frag_a QL1 ( .A1(J), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // jkffpc

`endif

`ifdef jkff
`else
`define jkff
module jkff( CLK , J, K, Q );
input CLK /* synthesis syn_isclock=1 */;
input J, K;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(CLK), .QD(N_1), .QR(GND), .QS(GND), .QZ(Q) );
frag_m I_2 ( .B1(Q), .B2(GND), .C1(GND), .C2(VCC), .D1(VCC), .D2(GND), .E1(VCC),
          .E2(Q), .NS(N_3), .OS(N_2), .OZ(N_1) );
frag_f I_1 ( .F1(K), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_3) );
frag_a QL1 ( .A1(J), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // jkff

`endif

`ifdef dffsc
`else
`define dffsc
module dffsc( CLK , CLR, D, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
wire N_3;
supply0 GND;

frag_f I_3 ( .F1(VCC), .F2(CLR), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_a I_2 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_q I_1 ( .QC(CLK), .QD(N_3), .QR(GND), .QS(GND), .QZ(Q) );
frag_m QL1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(GND), .D2(VCC), .E1(D),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(N_3) );

endmodule // dffsc

`endif

`ifdef dffpc
`else
`define dffpc
module dffpc( CLK , CLR, D, PRE, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input PRE /* synthesis syn_isclock=1 */;
input D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
wire N_3;
supply0 GND;

frag_f I_3 ( .F1(VCC), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_a I_2 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_q I_1 ( .QC(CLK), .QD(N_3), .QR(CLR), .QS(PRE), .QZ(Q) );
frag_m QL1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(D),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(N_3) );

endmodule // dffpc

`endif

`ifdef dffp
`else
`define dffp
module dffp( CLK , D, PRE, Q );
input CLK /* synthesis syn_isclock=1 */;
input PRE /* synthesis syn_isclock=1 */;
input D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
wire N_3;
supply0 GND;

frag_f I_3 ( .F1(VCC), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_a I_2 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_q I_1 ( .QC(CLK), .QD(N_3), .QR(GND), .QS(PRE), .QZ(Q) );
frag_m QL1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(D),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(N_3) );

endmodule // dffp

`endif

`ifdef dffepc
`else
`define dffepc
module dffepc( CLK , CLR, D, EN, PRE, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input PRE /* synthesis syn_isclock=1 */;
input D, EN;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply1 VCC;
supply0 GND;

frag_a I_3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_1) );
frag_m I_2 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(Q), .D2(GND), .E1(D),
          .E2(GND), .NS(N_3), .OS(N_1), .OZ(N_2) );
frag_q I_1 ( .QC(CLK), .QD(N_2), .QR(CLR), .QS(PRE), .QZ(Q) );
frag_f QL1 ( .F1(EN), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_3) );

endmodule // dffepc

`endif

`ifdef dffe
`else
`define dffe
module dffe( CLK , D, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input D, EN;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply1 VCC;
supply0 GND;

frag_a I_3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_1) );
frag_m I_2 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(Q), .D2(GND), .E1(D),
          .E2(GND), .NS(N_3), .OS(N_1), .OZ(N_2) );
frag_q I_1 ( .QC(CLK), .QD(N_2), .QR(GND), .QS(GND), .QZ(Q) );
frag_f QL1 ( .F1(EN), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_3) );

endmodule // dffe

`endif

`ifdef dffc
`else
`define dffc
module dffc( CLK , CLR, D, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
wire N_3;
supply0 GND;

frag_f I_3 ( .F1(VCC), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_a I_2 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_q I_1 ( .QC(CLK), .QD(N_3), .QR(CLR), .QS(GND), .QZ(Q) );
frag_m QL1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(D),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(N_3) );

endmodule // dffc

`endif

`ifdef dff
`else
`define dff
module dff( CLK , D, Q );
input CLK /* synthesis syn_isclock=1 */;
input D;
output Q;
parameter ql_gate = `LOGIC;
supply0 GND;
wire N_1;
supply1 VCC;
wire N_2;
wire N_3;

frag_m I_3 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(GND), .E1(D),
          .E2(GND), .NS(N_2), .OS(N_3), .OZ(N_1) );
frag_q I_2 ( .QC(CLK), .QD(N_1), .QR(GND), .QS(GND), .QZ(Q) );
frag_a I_1 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_3) );
frag_f QL1 ( .F1(VCC), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );

endmodule // dff

`endif

`ifdef udcnt6
`else
`define udcnt6
module udcnt6( CLK , CLR, ENP, ENT, UP, Q, RCO );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input ENP, ENT;
 output [5:0] Q;
output RCO;
input UP;
wire N_1;
wire N_2;

udcnt3b I_2 ( .CLK(CLK), .CLR(CLR), .ENP(N_2), .ENT(ENP), .Q({ Q[3],Q[4],Q[5] }),
           .RCO(N_1), .UP(UP) );
udcnt3a I_3 ( .CLK(CLK), .CLR(CLR), .ENP(ENP), .ENT(ENT), .Q({ Q[0],Q[1],Q[2] }),
           .RCO(N_2), .UP(UP) );
nand2i1 I_1 ( .A(N_2), .B(N_1), .Q(RCO) );

endmodule // udcnt6

`endif

`ifdef udcnt3
`else
`define udcnt3
module udcnt3( CLK , CLR, ENP, ENT, UP, Q, RCO );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input ENP, ENT;
 output [2:0] Q;
output RCO;
input UP;

udcnt3a I_1 ( .CLK(CLK), .CLR(CLR), .ENP(ENP), .ENT(ENT), .Q({ Q[0],Q[1],Q[2] }),
           .RCO(RCO), .UP(UP) );

endmodule // udcnt3

`endif

`ifdef udcnt12
`else
`define udcnt12
module udcnt12( CLK , CLR, ENP, ENT, UP, Q, RCO );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input ENP, ENT;
 output [11:0] Q;
output RCO;
input UP;
wire N_1;
wire N_2;
wire N_3;
wire N_4;

udcnt3b I_2 ( .CLK(CLK), .CLR(CLR), .ENP(N_4), .ENT(N_2), .Q({ Q[9],Q[10],Q[11] }),
           .RCO(N_1), .UP(UP) );
udcnt3b I_3 ( .CLK(CLK), .CLR(CLR), .ENP(N_4), .ENT(N_3), .Q({ Q[6],Q[7],Q[8] }),
           .RCO(N_2), .UP(UP) );
udcnt3b I_4 ( .CLK(CLK), .CLR(CLR), .ENP(N_4), .ENT(ENP), .Q({ Q[3],Q[4],Q[5] }),
           .RCO(N_3), .UP(UP) );
udcnt3a I_5 ( .CLK(CLK), .CLR(CLR), .ENP(ENP), .ENT(ENT), .Q({ Q[0],Q[1],Q[2] }),
           .RCO(N_4), .UP(UP) );
nand2i1 I_1 ( .A(N_4), .B(N_1), .Q(RCO) );

endmodule // udcnt12

`endif

`ifdef ucntx8
`else
`define ucntx8
module ucntx8( CLK , CLR, D, EN, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [7:0] D;
input EN, LOAD;
 output [7:0] Q;
wire N_1;
wire N_2;

uctxcar1 I_1 ( .ACO1(N_2), .CLK(CLK), .CLR(CLR), .D({ D[0],D[1] }), .ENG(EN),
            .LOAD(LOAD), .Q({ Q[0],Q[1] }) );
ucntx4c I_2 ( .CLK(CLK), .CLR(CLR), .D({ D[4],D[5],D[6],D[7] }), .ENG(EN), .ENP(N_2), .ENT(N_1),
           .LOAD(LOAD), .Q({ Q[4],Q[5],Q[6],Q[7] }) );
ucntx4a I_3 ( .CLK(CLK), .CLR(CLR), .D({ D[0],D[1],D[2],D[3] }), .ENG(EN), .LOAD(LOAD),
           .Q({ Q[0],Q[1],Q[2],Q[3] }), .RCO(N_1) );

endmodule // ucntx8

`endif

`ifdef ucntx4
`else
`define ucntx4
module ucntx4( CLK , CLR, D, EN, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [3:0] D;
input EN, LOAD;
 output [3:0] Q;
supply0 GND;

ucntx4c I_1 ( .CLK(CLK), .CLR(CLR), .D({ D[0],D[1],D[2],D[3] }), .ENG(EN), .ENP(GND), .ENT(GND),
           .LOAD(LOAD), .Q({ Q[0],Q[1],Q[2],Q[3] }) );

endmodule // ucntx4

`endif

`ifdef ucntx32
`else
`define ucntx32
module ucntx32( CLK , CLR, D, EN, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [31:0] D;
input EN, LOAD;
 output [31:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;

ucntx4c I_1 ( .CLK(CLK), .CLR(CLR), .D({ D[28],D[29],D[30],D[31] }), .ENG(EN), .ENP(N_14),
           .ENT(N_11), .LOAD(LOAD), .Q({ Q[28],Q[29],Q[30],Q[31] }) );
ucntx4a I_2 ( .CLK(CLK), .CLR(CLR), .D({ D[0],D[1],D[2],D[3] }), .ENG(EN), .LOAD(LOAD),
           .Q({ Q[0],Q[1],Q[2],Q[3] }), .RCO(N_1) );
ucntx4b I_3 ( .CLK(CLK), .CLR(CLR), .D({ D[16],D[17],D[18],D[19] }), .ENG(EN), .ENP(N_9),
           .ENT(N_8), .LOAD(LOAD), .Q({ Q[16],Q[17],Q[18],Q[19] }), .RCO(N_7) );
ucntx4b I_4 ( .CLK(CLK), .CLR(CLR), .D({ D[20],D[21],D[22],D[23] }), .ENG(EN), .ENP(N_10),
           .ENT(N_7), .LOAD(LOAD), .Q({ Q[20],Q[21],Q[22],Q[23] }), .RCO(N_12) );
ucntx4b I_5 ( .CLK(CLK), .CLR(CLR), .D({ D[24],D[25],D[26],D[27] }), .ENG(EN), .ENP(N_13),
           .ENT(N_12), .LOAD(LOAD), .Q({ Q[24],Q[25],Q[26],Q[27] }), .RCO(N_11) );
ucntx4b I_6 ( .CLK(CLK), .CLR(CLR), .D({ D[12],D[13],D[14],D[15] }), .ENG(EN), .ENP(N_6),
           .ENT(N_2), .LOAD(LOAD), .Q({ Q[12],Q[13],Q[14],Q[15] }), .RCO(N_8) );
ucntx4b I_7 ( .CLK(CLK), .CLR(CLR), .D({ D[8],D[9],D[10],D[11] }), .ENG(EN), .ENP(N_5),
           .ENT(N_3), .LOAD(LOAD), .Q({ Q[8],Q[9],Q[10],Q[11] }), .RCO(N_2) );
ucntx4b I_8 ( .CLK(CLK), .CLR(CLR), .D({ D[4],D[5],D[6],D[7] }), .ENG(EN), .ENP(N_4), .ENT(N_1),
           .LOAD(LOAD), .Q({ Q[4],Q[5],Q[6],Q[7] }), .RCO(N_3) );
uctxcar2 I_9 ( .ACO1(N_13), .ACO2(N_14), .CLK(CLK), .CLR(CLR), .D({ D[0],D[1] }),
            .ENG(EN), .LOAD(LOAD) );
uctxcar2 I_10 ( .ACO1(N_9), .ACO2(N_10), .CLK(CLK), .CLR(CLR), .D({ D[0],D[1] }),
             .ENG(EN), .LOAD(LOAD) );
uctxcar3 I_11 ( .ACO1(N_4), .ACO2(N_5), .ACO3(N_6), .CLK(CLK), .CLR(CLR),
             .D({ D[0],D[1] }), .ENG(EN), .LOAD(LOAD), .Q({ Q[0],Q[1] }) );

endmodule // ucntx32

`endif

`ifdef ucntx24
`else
`define ucntx24
module ucntx24( CLK , CLR, D, EN, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [23:0] D;
input EN, LOAD;
 output [23:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;

uctxcar3 I_1 ( .ACO1(N_4), .ACO2(N_5), .ACO3(N_6), .CLK(CLK), .CLR(CLR),
            .D({ D[0],D[1] }), .ENG(EN), .LOAD(LOAD), .Q({ Q[0],Q[1] }) );
uctxcar2 I_2 ( .ACO1(N_9), .ACO2(N_10), .CLK(CLK), .CLR(CLR), .D({ D[0],D[1] }),
            .ENG(EN), .LOAD(LOAD) );
ucntx4c I_3 ( .CLK(CLK), .CLR(CLR), .D({ D[20],D[21],D[22],D[23] }), .ENG(EN), .ENP(N_10),
           .ENT(N_8), .LOAD(LOAD), .Q({ Q[20],Q[21],Q[22],Q[23] }) );
ucntx4b I_4 ( .CLK(CLK), .CLR(CLR), .D({ D[16],D[17],D[18],D[19] }), .ENG(EN), .ENP(N_9),
           .ENT(N_7), .LOAD(LOAD), .Q({ Q[16],Q[17],Q[18],Q[19] }), .RCO(N_8) );
ucntx4b I_5 ( .CLK(CLK), .CLR(CLR), .D({ D[12],D[13],D[14],D[15] }), .ENG(EN), .ENP(N_6),
           .ENT(N_2), .LOAD(LOAD), .Q({ Q[12],Q[13],Q[14],Q[15] }), .RCO(N_7) );
ucntx4b I_6 ( .CLK(CLK), .CLR(CLR), .D({ D[8],D[9],D[10],D[11] }), .ENG(EN), .ENP(N_5),
           .ENT(N_3), .LOAD(LOAD), .Q({ Q[8],Q[9],Q[10],Q[11] }), .RCO(N_2) );
ucntx4b I_7 ( .CLK(CLK), .CLR(CLR), .D({ D[4],D[5],D[6],D[7] }), .ENG(EN), .ENP(N_4), .ENT(N_1),
           .LOAD(LOAD), .Q({ Q[4],Q[5],Q[6],Q[7] }), .RCO(N_3) );
ucntx4a I_8 ( .CLK(CLK), .CLR(CLR), .D({ D[0],D[1],D[2],D[3] }), .ENG(EN), .LOAD(LOAD),
           .Q({ Q[0],Q[1],Q[2],Q[3] }), .RCO(N_1) );

endmodule // ucntx24

`endif

`ifdef ucntx16
`else
`define ucntx16
module ucntx16( CLK , CLR, D, EN, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [15:0] D;
input EN, LOAD;
 output [15:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;

ucntx4c I_1 ( .CLK(CLK), .CLR(CLR), .D({ D[12],D[13],D[14],D[15] }), .ENG(EN), .ENP(N_6),
           .ENT(N_2), .LOAD(LOAD), .Q({ Q[12],Q[13],Q[14],Q[15] }) );
uctxcar3 I_2 ( .ACO1(N_4), .ACO2(N_5), .ACO3(N_6), .CLK(CLK), .CLR(CLR),
            .D({ D[0],D[1] }), .ENG(EN), .LOAD(LOAD), .Q({ Q[0],Q[1] }) );
ucntx4b I_3 ( .CLK(CLK), .CLR(CLR), .D({ D[8],D[9],D[10],D[11] }), .ENG(EN), .ENP(N_5),
           .ENT(N_3), .LOAD(LOAD), .Q({ Q[8],Q[9],Q[10],Q[11] }), .RCO(N_2) );
ucntx4b I_4 ( .CLK(CLK), .CLR(CLR), .D({ D[4],D[5],D[6],D[7] }), .ENG(EN), .ENP(N_4), .ENT(N_1),
           .LOAD(LOAD), .Q({ Q[4],Q[5],Q[6],Q[7] }), .RCO(N_3) );
ucntx4a I_5 ( .CLK(CLK), .CLR(CLR), .D({ D[0],D[1],D[2],D[3] }), .ENG(EN), .LOAD(LOAD),
           .Q({ Q[0],Q[1],Q[2],Q[3] }), .RCO(N_1) );

endmodule // ucntx16

`endif

`ifdef ucntl8
`else
`define ucntl8
module ucntl8( CLK , CLR, D, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [7:0] D;
input LOAD;
 output [7:0] Q;
wire N_1;
supply0 GND;

uctlcar1 I_1 ( .ACO1(N_1), .CLK(CLK), .CLR(CLR), .D({ D[0],D[1],D[2],D[3] }), .LOAD(LOAD),
            .Q({ Q[0],Q[1],Q[2],Q[3] }) );
ucntl4c I_2 ( .CLK(CLK), .CLR(CLR), .D({ D[4],D[5],D[6],D[7] }), .ENP(N_1), .ENT(GND),
           .LOAD(LOAD), .Q({ Q[4],Q[5],Q[6],Q[7] }) );
ucntl4c I_3 ( .CLK(CLK), .CLR(CLR), .D({ D[0],D[1],D[2],D[3] }), .ENP(GND), .ENT(GND),
           .LOAD(LOAD), .Q({ Q[0],Q[1],Q[2],Q[3] }) );

endmodule // ucntl8

`endif

`ifdef ucntl4
`else
`define ucntl4
module ucntl4( CLK , CLR, D, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [3:0] D;
input LOAD;
 output [3:0] Q;
supply0 GND;

ucntl4c I_1 ( .CLK(CLK), .CLR(CLR), .D({ D[0],D[1],D[2],D[3] }), .ENP(GND), .ENT(GND),
           .LOAD(LOAD), .Q({ Q[0],Q[1],Q[2],Q[3] }) );

endmodule // ucntl4

`endif

`ifdef ucntl32
`else
`define ucntl32
module ucntl32( CLK , CLR, D, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [31:0] D;
input LOAD;
 output [31:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;

uctlcar3 I_1 ( .ACO1(N_8), .ACO2(N_11), .ACO3(N_14), .CLK(CLK), .CLR(CLR),
            .D({ D[0],D[1] }), .LOAD(LOAD) );
uctlcar2 I_2 ( .ACO1(N_9), .ACO2(N_12), .CLK(CLK), .CLR(CLR), .D({ D[0],D[1] }),
            .LOAD(LOAD) );
uctlcar2 I_3 ( .ACO1(N_10), .ACO2(N_13), .CLK(CLK), .CLR(CLR), .D({ D[0],D[1] }),
            .LOAD(LOAD) );
ucntl4b I_4 ( .CLK(CLK), .CLR(CLR), .D({ D[24],D[25],D[26],D[27] }), .ENP(N_11), .ENT(N_3),
           .LOAD(LOAD), .Q({ Q[24],Q[25],Q[26],Q[27] }), .RCO(N_2) );
ucntl4b I_5 ( .CLK(CLK), .CLR(CLR), .D({ D[20],D[21],D[22],D[23] }), .ENP(N_8), .ENT(N_4),
           .LOAD(LOAD), .Q({ Q[20],Q[21],Q[22],Q[23] }), .RCO(N_3) );
ucntl4b I_6 ( .CLK(CLK), .CLR(CLR), .D({ D[16],D[17],D[18],D[19] }), .ENP(N_12), .ENT(N_5),
           .LOAD(LOAD), .Q({ Q[16],Q[17],Q[18],Q[19] }), .RCO(N_4) );
ucntl4b I_7 ( .CLK(CLK), .CLR(CLR), .D({ D[12],D[13],D[14],D[15] }), .ENP(N_9), .ENT(N_6),
           .LOAD(LOAD), .Q({ Q[12],Q[13],Q[14],Q[15] }), .RCO(N_5) );
ucntl4b I_8 ( .CLK(CLK), .CLR(CLR), .D({ D[8],D[9],D[10],D[11] }), .ENP(N_13), .ENT(N_7),
           .LOAD(LOAD), .Q({ Q[8],Q[9],Q[10],Q[11] }), .RCO(N_6) );
ucntl4b I_9 ( .CLK(CLK), .CLR(CLR), .D({ D[4],D[5],D[6],D[7] }), .ENP(N_10), .ENT(N_1),
           .LOAD(LOAD), .Q({ Q[4],Q[5],Q[6],Q[7] }), .RCO(N_7) );
ucntl4a I_10 ( .CLK(CLK), .CLR(CLR), .D({ D[0],D[1],D[2],D[3] }), .LOAD(LOAD), .Q({ Q[0],Q[1],Q[2],Q[3] }),
            .RCO(N_1) );
ucntl4c I_11 ( .CLK(CLK), .CLR(CLR), .D({ D[28],D[29],D[30],D[31] }), .ENP(N_14), .ENT(N_2),
            .LOAD(LOAD), .Q({ Q[28],Q[29],Q[30],Q[31] }) );

endmodule // ucntl32

`endif

`ifdef ucntl24
`else
`define ucntl24
module ucntl24( CLK , CLR, D, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [23:0] D;
input LOAD;
 output [23:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;

uctlcar2 I_1 ( .ACO1(N_4), .ACO2(N_5), .CLK(CLK), .CLR(CLR), .D({ D[0],D[1] }),
            .LOAD(LOAD) );
uctlcar3 I_2 ( .ACO1(N_8), .ACO2(N_9), .ACO3(N_10), .CLK(CLK), .CLR(CLR),
            .D({ D[0],D[1] }), .LOAD(LOAD) );
ucntl4b I_3 ( .CLK(CLK), .CLR(CLR), .D({ D[16],D[17],D[18],D[19] }), .ENP(N_9), .ENT(N_7),
           .LOAD(LOAD), .Q({ Q[16],Q[17],Q[18],Q[19] }), .RCO(N_6) );
ucntl4b I_4 ( .CLK(CLK), .CLR(CLR), .D({ D[12],D[13],D[14],D[15] }), .ENP(N_8), .ENT(N_2),
           .LOAD(LOAD), .Q({ Q[12],Q[13],Q[14],Q[15] }), .RCO(N_7) );
ucntl4b I_5 ( .CLK(CLK), .CLR(CLR), .D({ D[8],D[9],D[10],D[11] }), .ENP(N_5), .ENT(N_3),
           .LOAD(LOAD), .Q({ Q[8],Q[9],Q[10],Q[11] }), .RCO(N_2) );
ucntl4b I_6 ( .CLK(CLK), .CLR(CLR), .D({ D[4],D[5],D[6],D[7] }), .ENP(N_4), .ENT(N_1),
           .LOAD(LOAD), .Q({ Q[4],Q[5],Q[6],Q[7] }), .RCO(N_3) );
ucntl4a I_7 ( .CLK(CLK), .CLR(CLR), .D({ D[0],D[1],D[2],D[3] }), .LOAD(LOAD), .Q({ Q[0],Q[1],Q[2],Q[3] }),
           .RCO(N_1) );
ucntl4c I_8 ( .CLK(CLK), .CLR(CLR), .D({ D[20],D[21],D[22],D[23] }), .ENP(N_10), .ENT(N_6),
           .LOAD(LOAD), .Q({ Q[20],Q[21],Q[22],Q[23] }) );

endmodule // ucntl24

`endif

`ifdef ucntl16
`else
`define ucntl16
module ucntl16( CLK , CLR, D, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [15:0] D;
input LOAD;
 output [15:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;

ucntl4c I_1 ( .CLK(CLK), .CLR(CLR), .D({ D[12],D[13],D[14],D[15] }), .ENP(N_6), .ENT(N_2),
           .LOAD(LOAD), .Q({ Q[12],Q[13],Q[14],Q[15] }) );
uctlcar3 I_2 ( .ACO1(N_4), .ACO2(N_5), .ACO3(N_6), .CLK(CLK), .CLR(CLR),
            .D({ D[0],D[1] }), .LOAD(LOAD) );
ucntl4b I_3 ( .CLK(CLK), .CLR(CLR), .D({ D[8],D[9],D[10],D[11] }), .ENP(N_5), .ENT(N_3),
           .LOAD(LOAD), .Q({ Q[8],Q[9],Q[10],Q[11] }), .RCO(N_2) );
ucntl4b I_4 ( .CLK(CLK), .CLR(CLR), .D({ D[4],D[5],D[6],D[7] }), .ENP(N_4), .ENT(N_1),
           .LOAD(LOAD), .Q({ Q[4],Q[5],Q[6],Q[7] }), .RCO(N_3) );
ucntl4a I_5 ( .CLK(CLK), .CLR(CLR), .D({ D[0],D[1],D[2],D[3] }), .LOAD(LOAD), .Q({ Q[0],Q[1],Q[2],Q[3] }),
           .RCO(N_1) );

endmodule // ucntl16

`endif

`ifdef ucnte8
`else
`define ucnte8
module ucnte8( CLK , CLR, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input EN;
 output [7:0] Q;
wire N_1;
supply0 GND;

uctecar1 I_1 ( .ACO1(N_1), .CLK(CLK), .CLR(CLR), .ENG(EN), .Q({ Q[0],Q[1],Q[2],Q[3] }) );
ucnte4c I_2 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_1), .ENT(GND), .Q({ Q[4],Q[5],Q[6],Q[7] }) );
ucnte4c I_3 ( .CLK(CLK), .CLR(CLR), .ENG(GND), .ENP(EN), .ENT(GND), .Q({ Q[0],Q[1],Q[2],Q[3] }) );

endmodule // ucnte8

`endif

`ifdef ucnte4
`else
`define ucnte4
module ucnte4( CLK , CLR, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input EN;
 output [3:0] Q;
supply0 GND;

ucnte4c I_1 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(GND), .ENT(GND), .Q({ Q[0],Q[1],Q[2],Q[3] }) );

endmodule // ucnte4

`endif

`ifdef ucnte32
`else
`define ucnte32
module ucnte32( CLK , CLR, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input EN;
 output [31:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;

ucnte4b I_1 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_3), .ENT(N_13),
           .Q({ Q[24],Q[25],Q[26],Q[27] }), .RCO(N_14) );
ucnte4b I_2 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_2), .ENT(N_1),
           .Q({ Q[20],Q[21],Q[22],Q[23] }), .RCO(N_13) );
ucnte4b I_3 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_5), .ENT(N_6),
           .Q({ Q[16],Q[17],Q[18],Q[19] }), .RCO(N_1) );
ucnte4b I_4 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_10), .ENT(N_7),
           .Q({ Q[12],Q[13],Q[14],Q[15] }), .RCO(N_6) );
ucnte4b I_5 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_12), .ENT(N_8),
           .Q({ Q[8],Q[9],Q[10],Q[11] }), .RCO(N_7) );
ucnte4b I_6 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_11), .ENT(N_9),
           .Q({ Q[4],Q[5],Q[6],Q[7] }), .RCO(N_8) );
ucnte4a I_7 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .Q({ Q[0],Q[1],Q[2],Q[3] }), .RCO(N_9) );
ucnte4c I_8 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_4), .ENT(N_14),
           .Q({ Q[28],Q[29],Q[30],Q[31] }) );
upfecar2 QL9 ( .ACO1(N_10), .ACO2(N_5), .CLK(CLK), .CLR(CLR), .ENG(EN) );
upfecar2 QL10 ( .ACO1(N_11), .ACO2(N_12), .CLK(CLK), .CLR(CLR), .ENG(EN) );
upfecar3 QL11 ( .ACO1(N_2), .ACO2(N_3), .ACO3(N_4), .CLK(CLK), .CLR(CLR), .ENG(EN) );

endmodule // ucnte32

`endif

`ifdef ucnte24
`else
`define ucnte24
module ucnte24( CLK , CLR, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input EN;
 output [23:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;

ucnte4c I_1 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_6), .ENT(N_9),
           .Q({ Q[20],Q[21],Q[22],Q[23] }) );
ucnte4b I_2 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_7), .ENT(N_10),
           .Q({ Q[16],Q[17],Q[18],Q[19] }), .RCO(N_9) );
ucnte4b I_3 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_8), .ENT(N_1),
           .Q({ Q[12],Q[13],Q[14],Q[15] }), .RCO(N_10) );
ucnte4b I_4 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_5), .ENT(N_2),
           .Q({ Q[8],Q[9],Q[10],Q[11] }), .RCO(N_1) );
ucnte4b I_5 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_4), .ENT(N_3), .Q({ Q[4],Q[5],Q[6],Q[7] }),
           .RCO(N_2) );
ucnte4a I_6 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .Q({ Q[0],Q[1],Q[2],Q[3] }), .RCO(N_3) );
upfecar2 QL7 ( .ACO1(N_4), .ACO2(N_5), .CLK(CLK), .CLR(CLR), .ENG(EN) );
upfecar3 QL8 ( .ACO1(N_8), .ACO2(N_7), .ACO3(N_6), .CLK(CLK), .CLR(CLR), .ENG(EN) );

endmodule // ucnte24

`endif

`ifdef ucnte16
`else
`define ucnte16
module ucnte16( CLK , CLR, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input EN;
 output [15:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;

ucnte4c I_1 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_4), .ENT(N_2),
           .Q({ Q[12],Q[13],Q[14],Q[15] }) );
ucnte4b I_2 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_5), .ENT(N_3),
           .Q({ Q[8],Q[9],Q[10],Q[11] }), .RCO(N_2) );
ucnte4b I_3 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_6), .ENT(N_1), .Q({ Q[4],Q[5],Q[6],Q[7] }),
           .RCO(N_3) );
ucnte4a I_4 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .Q({ Q[0],Q[1],Q[2],Q[3] }), .RCO(N_1) );
upfecar3 QL5 ( .ACO1(N_6), .ACO2(N_5), .ACO3(N_4), .CLK(CLK), .CLR(CLR), .ENG(EN) );

endmodule // ucnte16

`endif

`ifdef rcnt8
`else
`define rcnt8
module rcnt8( CI , CLK, CLR, D, LOAD, CO, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input CI;
output CO;
 input [7:0] D;
input LOAD;
 output [7:0] Q;
wire N_1;

rcnt4 QL4 ( .CI(CI), .CLK(CLK), .CLR(CLR), .CO(N_1), .D({ D[3:0] }), .LOAD(LOAD),
         .Q({ Q[3:0] }) );
rcnt4 QL3 ( .CI(N_1), .CLK(CLK), .CLR(CLR), .CO(CO), .D({ D[7:4] }), .LOAD(LOAD),
         .Q({ Q[7:4] }) );

endmodule // rcnt8

`endif

`ifdef rcnt4
`else
`define rcnt4
module rcnt4( CI , CLK, CLR, D, LOAD, CO, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input CI;
output CO;
 input [3:0] D;
input LOAD;
 output [3:0] Q;
wire N_1;
supply1 VCC;
wire N_2;
wire N_3;
wire N_4;

and2i0 I_1 ( .A(N_1), .B(Q[3]), .Q(CO) );
ripbit QL1 ( .CI(N_3), .CLK(CLK), .CLR(CLR), .CO(N_1), .CX(Q[2]), .D(D[3]),
          .LOAD(LOAD), .Q(Q[3]) );
ripbit QL2 ( .CI(N_2), .CLK(CLK), .CLR(CLR), .CO(N_3), .CX(Q[1]), .D(D[2]),
          .LOAD(LOAD), .Q(Q[2]) );
ripbit QL3 ( .CI(N_4), .CLK(CLK), .CLR(CLR), .CO(N_2), .CX(Q[0]), .D(D[1]),
          .LOAD(LOAD), .Q(Q[1]) );
ripbit QL4 ( .CI(CI), .CLK(CLK), .CLR(CLR), .CO(N_4), .CX(VCC), .D(D[0]),
          .LOAD(LOAD), .Q(Q[0]) );

endmodule // rcnt4

`endif

`ifdef rcnt16
`else
`define rcnt16
module rcnt16( CI , CLK, CLR, D, LOAD, CO, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input CI;
output CO;
 input [15:0] D;
input LOAD;
 output [15:0] Q;
wire N_1;
wire N_2;
wire N_3;

rcnt4 QL8 ( .CI(CI), .CLK(CLK), .CLR(CLR), .CO(N_3), .D({ D[3:0] }), .LOAD(LOAD),
         .Q({ Q[3:0] }) );
rcnt4 QL7 ( .CI(N_3), .CLK(CLK), .CLR(CLR), .CO(N_2), .D({ D[7:4] }), .LOAD(LOAD),
         .Q({ Q[7:4] }) );
rcnt4 QL6 ( .CI(N_2), .CLK(CLK), .CLR(CLR), .CO(N_1), .D({ D[11:8] }), .LOAD(LOAD),
         .Q({ Q[11:8] }) );
rcnt4 QL5 ( .CI(N_1), .CLK(CLK), .CLR(CLR), .CO(CO), .D({ D[15:12] }), .LOAD(LOAD),
         .Q({ Q[15:12] }) );

endmodule // rcnt16

`endif

`ifdef dcntx8
`else
`define dcntx8
module dcntx8( CLK , CLR, D, EN, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [7:0] D;
input EN, LOAD;
 output [7:0] Q;
wire N_1;
wire N_2;

dctxcar1 I_1 ( .ACO1(N_2), .CLK(CLK), .CLR(CLR), .D({ D[1:0] }), .ENG(EN),
            .LOAD(LOAD), .Q({ Q[1:0] }) );
dcntx4a I_2 ( .CLK(CLK), .CLR(CLR), .D({ D[3:0] }), .ENG(EN), .LOAD(LOAD),
           .Q({ Q[3:0] }), .RCO(N_1) );
dcntx4c I_3 ( .CLK(CLK), .CLR(CLR), .D({ D[7:4] }), .ENG(EN), .ENP(N_2), .ENT(N_1),
           .LOAD(LOAD), .Q({ Q[7:4] }) );

endmodule // dcntx8

`endif

`ifdef dcntx4
`else
`define dcntx4
module dcntx4( CLK , CLR, D, EN, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [3:0] D;
input EN, LOAD;
 output [3:0] Q;
supply1 VCC;

dcntx4c I_1 ( .CLK(CLK), .CLR(CLR), .D({ D[3:0] }), .ENG(EN), .ENP(VCC), .ENT(VCC),
           .LOAD(LOAD), .Q({ Q[3:0] }) );

endmodule // dcntx4

`endif

`ifdef dcntx32
`else
`define dcntx32
module dcntx32( CLK , CLR, D, EN, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [31:0] D;
input EN, LOAD;
 output [31:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;

dctxcar2 I_1 ( .ACO1(N_13), .ACO2(N_14), .CLK(CLK), .CLR(CLR), .D({ D[1:0] }),
            .ENG(EN), .LOAD(LOAD) );
dctxcar2 I_2 ( .ACO1(N_9), .ACO2(N_10), .CLK(CLK), .CLR(CLR), .D({ D[1:0] }),
            .ENG(EN), .LOAD(LOAD) );
dctxcar3 I_3 ( .ACO1(N_4), .ACO2(N_5), .ACO3(N_6), .CLK(CLK), .CLR(CLR),
            .D({ D[1:0] }), .ENG(EN), .LOAD(LOAD), .Q({ Q[1:0] }) );
dcntx4c I_4 ( .CLK(CLK), .CLR(CLR), .D({ D[31:28] }), .ENG(EN), .ENP(N_14),
           .ENT(N_11), .LOAD(LOAD), .Q({ Q[31:28] }) );
dcntx4b I_5 ( .CLK(CLK), .CLR(CLR), .D({ D[27:24] }), .ENG(EN), .ENP(N_13),
           .ENT(N_12), .LOAD(LOAD), .Q({ Q[27:24] }), .RCO(N_11) );
dcntx4b I_6 ( .CLK(CLK), .CLR(CLR), .D({ D[23:20] }), .ENG(EN), .ENP(N_10),
           .ENT(N_7), .LOAD(LOAD), .Q({ Q[23:20] }), .RCO(N_12) );
dcntx4b I_7 ( .CLK(CLK), .CLR(CLR), .D({ D[19:16] }), .ENG(EN), .ENP(N_9),
           .ENT(N_8), .LOAD(LOAD), .Q({ Q[19:16] }), .RCO(N_7) );
dcntx4b I_8 ( .CLK(CLK), .CLR(CLR), .D({ D[15:12] }), .ENG(EN), .ENP(N_6),
           .ENT(N_2), .LOAD(LOAD), .Q({ Q[15:12] }), .RCO(N_8) );
dcntx4b I_9 ( .CLK(CLK), .CLR(CLR), .D({ D[11:8] }), .ENG(EN), .ENP(N_5),
           .ENT(N_3), .LOAD(LOAD), .Q({ Q[11:8] }), .RCO(N_2) );
dcntx4b I_10 ( .CLK(CLK), .CLR(CLR), .D({ D[7:4] }), .ENG(EN), .ENP(N_4),
            .ENT(N_1), .LOAD(LOAD), .Q({ Q[7:4] }), .RCO(N_3) );
dcntx4a I_11 ( .CLK(CLK), .CLR(CLR), .D({ D[3:0] }), .ENG(EN), .LOAD(LOAD),
            .Q({ Q[3:0] }), .RCO(N_1) );

endmodule // dcntx32

`endif

`ifdef dcntx24
`else
`define dcntx24
module dcntx24( CLK , CLR, D, EN, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [23:0] D;
input EN, LOAD;
 output [23:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;

dctxcar3 I_1 ( .ACO1(N_4), .ACO2(N_5), .ACO3(N_6), .CLK(CLK), .CLR(CLR),
            .D({ D[1:0] }), .ENG(EN), .LOAD(LOAD), .Q({ Q[1:0] }) );
dcntx4c I_2 ( .CLK(CLK), .CLR(CLR), .D({ D[23:20] }), .ENG(EN), .ENP(N_10),
           .ENT(N_8), .LOAD(LOAD), .Q({ Q[23:20] }) );
dcntx4b I_3 ( .CLK(CLK), .CLR(CLR), .D({ D[19:16] }), .ENG(EN), .ENP(N_9),
           .ENT(N_7), .LOAD(LOAD), .Q({ Q[19:16] }), .RCO(N_8) );
dcntx4b I_4 ( .CLK(CLK), .CLR(CLR), .D({ D[15:12] }), .ENG(EN), .ENP(N_6),
           .ENT(N_2), .LOAD(LOAD), .Q({ Q[15:12] }), .RCO(N_7) );
dcntx4b I_5 ( .CLK(CLK), .CLR(CLR), .D({ D[11:8] }), .ENG(EN), .ENP(N_5),
           .ENT(N_3), .LOAD(LOAD), .Q({ Q[11:8] }), .RCO(N_2) );
dcntx4b I_6 ( .CLK(CLK), .CLR(CLR), .D({ D[7:4] }), .ENG(EN), .ENP(N_4), .ENT(N_1),
           .LOAD(LOAD), .Q({ Q[7:4] }), .RCO(N_3) );
dcntx4a I_7 ( .CLK(CLK), .CLR(CLR), .D({ D[3:0] }), .ENG(EN), .LOAD(LOAD),
           .Q({ Q[3:0] }), .RCO(N_1) );
dctxcar2 I_8 ( .ACO1(N_9), .ACO2(N_10), .CLK(CLK), .CLR(CLR), .D({ D[1:0] }),
            .ENG(EN), .LOAD(LOAD) );

endmodule // dcntx24

`endif

`ifdef dcntx16
`else
`define dcntx16
module dcntx16( CLK , CLR, D, EN, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [15:0] D;
input EN, LOAD;
 output [15:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;

dcntx4c I_1 ( .CLK(CLK), .CLR(CLR), .D({ D[15:12] }), .ENG(EN), .ENP(N_6),
           .ENT(N_2), .LOAD(LOAD), .Q({ Q[15:12] }) );
dcntx4b I_2 ( .CLK(CLK), .CLR(CLR), .D({ D[11:8] }), .ENG(EN), .ENP(N_5),
           .ENT(N_3), .LOAD(LOAD), .Q({ Q[11:8] }), .RCO(N_2) );
dcntx4b I_3 ( .CLK(CLK), .CLR(CLR), .D({ D[7:4] }), .ENG(EN), .ENP(N_4), .ENT(N_1),
           .LOAD(LOAD), .Q({ Q[7:4] }), .RCO(N_3) );
dcntx4a I_4 ( .CLK(CLK), .CLR(CLR), .D({ D[3:0] }), .ENG(EN), .LOAD(LOAD),
           .Q({ Q[3:0] }), .RCO(N_1) );
dctxcar3 I_5 ( .ACO1(N_4), .ACO2(N_5), .ACO3(N_6), .CLK(CLK), .CLR(CLR),
            .D({ D[1:0] }), .ENG(EN), .LOAD(LOAD), .Q({ Q[1:0] }) );

endmodule // dcntx16

`endif

`ifdef dcntl8
`else
`define dcntl8
module dcntl8( CLK , CLR, D, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [7:0] D;
input LOAD;
 output [7:0] Q;
supply1 VCC;
wire N_1;

dctlcar1 I_1 ( .ACO1(N_1), .CLK(CLK), .CLR(CLR), .D({ D[3:0] }), .LOAD(LOAD),
            .Q({ Q[3:0] }) );
dcntl4c I_2 ( .CLK(CLK), .CLR(CLR), .D({ D[7:4] }), .ENP(N_1), .ENT(VCC),
           .LOAD(LOAD), .Q({ Q[7:4] }) );
dcntl4c I_3 ( .CLK(CLK), .CLR(CLR), .D({ D[3:0] }), .ENP(VCC), .ENT(VCC),
           .LOAD(LOAD), .Q({ Q[3:0] }) );

endmodule // dcntl8

`endif

`ifdef dcntl4
`else
`define dcntl4
module dcntl4( CLK , CLR, D, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [3:0] D;
input LOAD;
 output [3:0] Q;
supply1 VCC;

dcntl4c I_1 ( .CLK(CLK), .CLR(CLR), .D({ D[3:0] }), .ENP(VCC), .ENT(VCC),
           .LOAD(LOAD), .Q({ Q[3:0] }) );

endmodule // dcntl4

`endif

`ifdef dcntl32
`else
`define dcntl32
module dcntl32( CLK , CLR, D, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [31:0] D;
input LOAD;
 output [31:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;

dctlcar3 I_1 ( .ACO1(N_8), .ACO2(N_11), .ACO3(N_14), .CLK(CLK), .CLR(CLR),
            .D({ D[1:0] }), .LOAD(LOAD) );
dctlcar2 I_2 ( .ACO1(N_10), .ACO2(N_13), .CLK(CLK), .CLR(CLR), .D({ D[1:0] }),
            .LOAD(LOAD) );
dctlcar2 I_3 ( .ACO1(N_9), .ACO2(N_12), .CLK(CLK), .CLR(CLR), .D({ D[1:0] }),
            .LOAD(LOAD) );
dcntl4b I_4 ( .CLK(CLK), .CLR(CLR), .D({ D[27:24] }), .ENP(N_11), .ENT(N_3),
           .LOAD(LOAD), .Q({ Q[27:24] }), .RCO(N_2) );
dcntl4b I_5 ( .CLK(CLK), .CLR(CLR), .D({ D[23:20] }), .ENP(N_8), .ENT(N_4),
           .LOAD(LOAD), .Q({ Q[23:20] }), .RCO(N_3) );
dcntl4b I_6 ( .CLK(CLK), .CLR(CLR), .D({ D[19:16] }), .ENP(N_12), .ENT(N_5),
           .LOAD(LOAD), .Q({ Q[19:16] }), .RCO(N_4) );
dcntl4b I_7 ( .CLK(CLK), .CLR(CLR), .D({ D[15:12] }), .ENP(N_9), .ENT(N_6),
           .LOAD(LOAD), .Q({ Q[15:12] }), .RCO(N_5) );
dcntl4b I_8 ( .CLK(CLK), .CLR(CLR), .D({ D[11:8] }), .ENP(N_13), .ENT(N_7),
           .LOAD(LOAD), .Q({ Q[11:8] }), .RCO(N_6) );
dcntl4b I_9 ( .CLK(CLK), .CLR(CLR), .D({ D[7:4] }), .ENP(N_10), .ENT(N_1),
           .LOAD(LOAD), .Q({ Q[7:4] }), .RCO(N_7) );
dcntl4a I_10 ( .CLK(CLK), .CLR(CLR), .D({ D[3:0] }), .LOAD(LOAD), .Q({ Q[3:0] }),
            .RCO(N_1) );
dcntl4c I_11 ( .CLK(CLK), .CLR(CLR), .D({ D[31:28] }), .ENP(N_14), .ENT(N_2),
            .LOAD(LOAD), .Q({ Q[31:28] }) );

endmodule // dcntl32

`endif

`ifdef dcntl24
`else
`define dcntl24
module dcntl24( CLK , CLR, D, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [23:0] D;
input LOAD;
 output [23:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;

dcntl4c I_1 ( .CLK(CLK), .CLR(CLR), .D({ D[23:20] }), .ENP(N_10), .ENT(N_6),
           .LOAD(LOAD), .Q({ Q[23:20] }) );
dctlcar3 I_2 ( .ACO1(N_8), .ACO2(N_9), .ACO3(N_10), .CLK(CLK), .CLR(CLR),
            .D({ D[1:0] }), .LOAD(LOAD) );
dcntl4b I_3 ( .CLK(CLK), .CLR(CLR), .D({ D[19:16] }), .ENP(N_9), .ENT(N_7),
           .LOAD(LOAD), .Q({ Q[19:16] }), .RCO(N_6) );
dcntl4b I_4 ( .CLK(CLK), .CLR(CLR), .D({ D[15:12] }), .ENP(N_8), .ENT(N_2),
           .LOAD(LOAD), .Q({ Q[15:12] }), .RCO(N_7) );
dcntl4b I_5 ( .CLK(CLK), .CLR(CLR), .D({ D[11:8] }), .ENP(N_5), .ENT(N_3),
           .LOAD(LOAD), .Q({ Q[11:8] }), .RCO(N_2) );
dcntl4b I_6 ( .CLK(CLK), .CLR(CLR), .D({ D[7:4] }), .ENP(N_4), .ENT(N_1),
           .LOAD(LOAD), .Q({ Q[7:4] }), .RCO(N_3) );
dcntl4a I_7 ( .CLK(CLK), .CLR(CLR), .D({ D[3:0] }), .LOAD(LOAD), .Q({ Q[3:0] }),
           .RCO(N_1) );
dctlcar2 I_8 ( .ACO1(N_4), .ACO2(N_5), .CLK(CLK), .CLR(CLR), .D({ D[1:0] }),
            .LOAD(LOAD) );

endmodule // dcntl24

`endif

`ifdef dcntl16
`else
`define dcntl16
module dcntl16( CLK , CLR, D, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [15:0] D;
input LOAD;
 output [15:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;

dctlcar3 I_1 ( .ACO1(N_4), .ACO2(N_5), .ACO3(N_6), .CLK(CLK), .CLR(CLR),
            .D({ D[1:0] }), .LOAD(LOAD) );
dcntl4b I_2 ( .CLK(CLK), .CLR(CLR), .D({ D[11:8] }), .ENP(N_5), .ENT(N_3),
           .LOAD(LOAD), .Q({ Q[11:8] }), .RCO(N_2) );
dcntl4b I_3 ( .CLK(CLK), .CLR(CLR), .D({ D[7:4] }), .ENP(N_4), .ENT(N_1),
           .LOAD(LOAD), .Q({ Q[7:4] }), .RCO(N_3) );
dcntl4a I_4 ( .CLK(CLK), .CLR(CLR), .D({ D[3:0] }), .LOAD(LOAD), .Q({ Q[3:0] }),
           .RCO(N_1) );
dcntl4c I_5 ( .CLK(CLK), .CLR(CLR), .D({ D[15:12] }), .ENP(N_6), .ENT(N_2),
           .LOAD(LOAD), .Q({ Q[15:12] }) );

endmodule // dcntl16

`endif

`ifdef dcnte8
`else
`define dcnte8
module dcnte8( CLK , CLR, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input EN;
 output [7:0] Q;
wire N_1;
supply1 VCC;

dctecar1 I_1 ( .ACO1(N_1), .CLK(CLK), .CLR(CLR), .ENG(EN), .Q({ Q[3:0] }) );
dcnte4c I_2 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_1), .ENT(VCC), .Q({ Q[7:4] }) );
dcnte4c I_3 ( .CLK(CLK), .CLR(CLR), .ENG(VCC), .ENP(EN), .ENT(VCC), .Q({ Q[3:0] }) );

endmodule // dcnte8

`endif

`ifdef dcnte4
`else
`define dcnte4
module dcnte4( CLK , CLR, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input EN;
 output [3:0] Q;
supply1 VCC;

dcnte4c I_1 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(VCC), .ENT(VCC), .Q({ Q[3:0] }) );

endmodule // dcnte4

`endif

`ifdef dcnte32
`else
`define dcnte32
module dcnte32( CLK , CLR, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input EN;
 output [31:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;

dcnte4c I_1 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_4), .ENT(N_14),
           .Q({ Q[31:28] }) );
dcnte4b I_2 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_3), .ENT(N_13),
           .Q({ Q[27:24] }), .RCO(N_14) );
dcnte4b I_3 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_2), .ENT(N_1),
           .Q({ Q[23:20] }), .RCO(N_13) );
dcnte4b I_4 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_5), .ENT(N_6),
           .Q({ Q[19:16] }), .RCO(N_1) );
dcnte4b I_5 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_10), .ENT(N_7),
           .Q({ Q[15:12] }), .RCO(N_6) );
dcnte4b I_6 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_12), .ENT(N_8),
           .Q({ Q[11:8] }), .RCO(N_7) );
dcnte4b I_7 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_11), .ENT(N_9),
           .Q({ Q[7:4] }), .RCO(N_8) );
dcnte4a I_8 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .Q({ Q[3:0] }), .RCO(N_9) );
dnfecar3 QL9 ( .ACO1(N_2), .ACO2(N_3), .ACO3(N_4), .CLK(CLK), .CLR(CLR), .ENG(EN) );
dnfecar2 QL10 ( .ACO1(N_10), .ACO2(N_5), .CLK(CLK), .CLR(CLR), .ENG(EN) );
dnfecar2 QL11 ( .ACO1(N_11), .ACO2(N_12), .CLK(CLK), .CLR(CLR), .ENG(EN) );

endmodule // dcnte32

`endif

`ifdef dcnte24
`else
`define dcnte24
module dcnte24( CLK , CLR, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input EN;
 output [23:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;

dcnte4b I_4 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_7), .ENT(N_10),
           .Q({ Q[19:16] }), .RCO(N_9) );
dcnte4b I_5 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_8), .ENT(N_1),
           .Q({ Q[15:12] }), .RCO(N_10) );
dcnte4b I_6 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_5), .ENT(N_2),
           .Q({ Q[11:8] }), .RCO(N_1) );
dcnte4b I_7 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_4), .ENT(N_3), .Q({ Q[7:4] }),
           .RCO(N_2) );
dcnte4a I_8 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .Q({ Q[3:0] }), .RCO(N_3) );
dcnte4c I_9 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_6), .ENT(N_9),
           .Q({ Q[23:20] }) );
dnfecar2 QL2 ( .ACO1(N_4), .ACO2(N_5), .CLK(CLK), .CLR(CLR), .ENG(EN) );
dnfecar3 QL7 ( .ACO1(N_8), .ACO2(N_7), .ACO3(N_6), .CLK(CLK), .CLR(CLR), .ENG(EN) );

endmodule // dcnte24

`endif

`ifdef dcnte16
`else
`define dcnte16
module dcnte16( CLK , CLR, EN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input EN;
 output [15:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;

dcnte4c I_1 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_4), .ENT(N_2),
           .Q({ Q[15:12] }) );
dcnte4b I_2 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_5), .ENT(N_3),
           .Q({ Q[11:8] }), .RCO(N_2) );
dcnte4b I_3 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .ENP(N_6), .ENT(N_1), .Q({ Q[7:4] }),
           .RCO(N_3) );
dcnte4a I_4 ( .CLK(CLK), .CLR(CLR), .ENG(EN), .Q({ Q[3:0] }), .RCO(N_1) );
dnfecar3 QL5 ( .ACO1(N_6), .ACO2(N_5), .ACO3(N_4), .CLK(CLK), .CLR(CLR), .ENG(EN) );

endmodule // dcnte16

`endif

`ifdef and6i6
`else
`define and6i6
module and6i6( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(VCC), .A2(D), .A3(VCC), .A4(E), .A5(VCC), .A6(F), .AZ(N_2) );
frag_f I_1 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m QL3 ( .B1(GND), .B2(VCC), .C1(GND), .C2(VCC), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // and6i6

`endif

`ifdef and6i5
`else
`define and6i5
module and6i5( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(VCC), .A2(D), .A3(VCC), .A4(E), .A5(VCC), .A6(F), .AZ(N_2) );
frag_f I_1 ( .F1(A), .F2(GND), .F3(VCC), .F4(B), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m QL3 ( .B1(GND), .B2(VCC), .C1(GND), .C2(VCC), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // and6i5

`endif

`ifdef and6i4
`else
`define and6i4
module and6i4( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(A), .F2(D), .F3(B), .F4(E), .F5(VCC), .F6(F), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(C), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // and6i4

`endif

`ifdef and6i3
`else
`define and6i3
module and6i3( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;

frag_a QL1 ( .A1(A), .A2(D), .A3(B), .A4(E), .A5(C), .A6(F), .AZ(Q) );

endmodule // and6i3

`endif

`ifdef and6i2
`else
`define and6i2
module and6i2( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(A), .F2(GND), .F3(B), .F4(E), .F5(C), .F6(F), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(GND), .D2(VCC), .E1(D),
          .E2(GND), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // and6i2

`endif

`ifdef and6i1
`else
`define and6i1
module and6i1( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(D), .A2(GND), .A3(E), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(A), .F2(GND), .F3(B), .F4(GND), .F5(C), .F6(F), .FZ(N_1) );
frag_m QL3 ( .B1(GND), .B2(VCC), .C1(GND), .C2(VCC), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // and6i1

`endif

`ifdef and6i0
`else
`define and6i0
module and6i0( A , B, C, D, E, F, Q );
input A, B, C, D, E, F;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(D), .A2(GND), .A3(E), .A4(GND), .A5(F), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(A), .F2(GND), .F3(B), .F4(GND), .F5(C), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(GND), .B2(VCC), .C1(GND), .C2(VCC), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // and6i0

`endif

`ifdef and5i5
`else
`define and5i5
module and5i5( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(VCC), .A2(D), .A3(VCC), .A4(E), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(VCC), .F2(A), .F3(VCC), .F4(B), .F5(VCC), .F6(C), .FZ(N_1) );
frag_m QL3 ( .B1(GND), .B2(VCC), .C1(GND), .C2(VCC), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // and5i5

`endif

`ifdef and5i4
`else
`define and5i4
module and5i4( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(A), .F2(C), .F3(VCC), .F4(D), .F5(VCC), .F6(E), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(B), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // and5i4

`endif

`ifdef and5i3
`else
`define and5i3
module and5i3( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;

frag_a QL1 ( .A1(A), .A2(D), .A3(B), .A4(E), .A5(VCC), .A6(C), .AZ(Q) );

endmodule // and5i3

`endif

`ifdef and5i2
`else
`define and5i2
module and5i2( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
supply0 GND;

frag_a QL1 ( .A1(A), .A2(GND), .A3(B), .A4(D), .A5(C), .A6(E), .AZ(Q) );

endmodule // and5i2

`endif

`ifdef and5i1
`else
`define and5i1
module and5i1( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(A), .F2(GND), .F3(B), .F4(E), .F5(C), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(GND), .D2(VCC), .E1(D),
          .E2(GND), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // and5i1

`endif

`ifdef and5i0
`else
`define and5i0
module and5i0( A , B, C, D, E, Q );
input A, B, C, D, E;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(D), .A2(GND), .A3(E), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_f I_1 ( .F1(A), .F2(GND), .F3(B), .F4(GND), .F5(C), .F6(GND), .FZ(N_1) );
frag_m QL3 ( .B1(GND), .B2(VCC), .C1(GND), .C2(VCC), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // and5i0

`endif

`ifdef and4i4
`else
`define and4i4
module and4i4( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(VCC), .F2(B), .F3(VCC), .F4(C), .F5(VCC), .F6(D), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(A), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // and4i4

`endif

`ifdef and4i3
`else
`define and4i3
module and4i3( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;

frag_a QL1 ( .A1(A), .A2(D), .A3(VCC), .A4(B), .A5(VCC), .A6(C), .AZ(Q) );

endmodule // and4i3

`endif

`ifdef and4i2
`else
`define and4i2
module and4i2( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter syn_macro = 1, ql_pack = 1;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

frag_a QL1 ( .A1(A), .A2(GND), .A3(B), .A4(D), .A5(VCC), .A6(C), .AZ(Q) );

endmodule // and4i2

`endif

`ifdef and4i1
`else
`define and4i1
module and4i1( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
supply0 GND;

frag_a QL1 ( .A1(A), .A2(GND), .A3(B), .A4(GND), .A5(C), .A6(D), .AZ(Q) );

endmodule // and4i1

`endif

`ifdef and4i0
`else
`define and4i0
module and4i0( A , B, C, D, Q );
input A, B, C, D;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;
wire N_2;

frag_f I_2 ( .F1(A), .F2(GND), .F3(B), .F4(GND), .F5(C), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(GND), .D2(VCC), .E1(D),
          .E2(GND), .NS(N_1), .NZ(Q), .OS(N_2) );
frag_a QL3 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // and4i0

`endif

`ifdef and3i3
`else
`define and3i3
module and3i3( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;

frag_a QL1 ( .A1(VCC), .A2(A), .A3(VCC), .A4(B), .A5(VCC), .A6(C), .AZ(Q) );

endmodule // and3i3

`endif

`ifdef and3i2
`else
`define and3i2
module and3i2( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

frag_a QL1 ( .A1(A), .A2(GND), .A3(VCC), .A4(B), .A5(VCC), .A6(C), .AZ(Q) );

endmodule // and3i2

`endif

`ifdef and3i1
`else
`define and3i1
module and3i1( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

frag_a QL1 ( .A1(A), .A2(GND), .A3(B), .A4(GND), .A5(VCC), .A6(C), .AZ(Q) );

endmodule // and3i1

`endif

`ifdef and3i0
`else
`define and3i0
module and3i0( A , B, C, Q );
input A, B, C;
output Q;
parameter ql_gate = `LOGIC;
supply0 GND;

frag_a QL1 ( .A1(A), .A2(GND), .A3(B), .A4(GND), .A5(C), .A6(GND), .AZ(Q) );

endmodule // and3i0

`endif

`ifdef and2i2
`else
`define and2i2
module and2i2( A , B, Q );
input A, B;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

frag_a QL1 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(A), .A5(VCC), .A6(B), .AZ(Q) );

endmodule // and2i2

`endif

`ifdef and2i1
`else
`define and2i1
module and2i1( A , B, Q );
input A, B;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

frag_a QL1 ( .A1(A), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(B), .AZ(Q) );

endmodule // and2i1

`endif

`ifdef and2i0
`else
`define and2i0
module and2i0( A , B, Q );
input A, B;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

frag_a QL1 ( .A1(A), .A2(GND), .A3(B), .A4(GND), .A5(VCC), .A6(GND), .AZ(Q) );

endmodule // and2i0

`endif

`ifdef sub8
`else
`define sub8
module sub8( A , B, Q );
 input [7:0] A;
 input [7:0] B;
 output [7:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;
wire N_15;
wire N_16;
wire N_17;
wire N_18;
wire N_19;
wire N_20;
wire N_21;
wire N_22;
wire N_23;
wire N_24;
wire N_25;
wire N_26;
wire N_27;
supply0 GND;
wire N_28;

csamuxa QL1 ( .A(N_18), .Q(Q[6]), .S00(N_21), .S01(N_17), .S1(N_19) );
csamuxb QL2 ( .A(N_15), .B(N_16), .Q(Q[7]), .S00(N_21), .S01(N_17), .S1(N_19) );
csamuxc QL3 ( .A(N_26), .B(N_27), .Q(N_19), .S00(N_5), .S01(N_6), .S1(N_8) );
csamuxd QL4 ( .A(N_4), .Q(Q[3]), .S00(N_5), .S01(N_6), .S1(N_24) );
csamuxd QL5 ( .A(N_14), .Q(Q[5]), .S00(N_20), .S01(N_22), .S1(N_19) );
mux4x6 QL6 ( .A(N_28), .B(N_28), .C(N_28), .D(N_28), .Q(Q[1]), .S0(N_7), .S1(B[1]) );
muxb2dx2 QL7 ( .A(N_13), .B(N_12), .C(GND), .D(GND), .Q(N_21), .S(N_10), .T(N_20) );
muxc2dx2 QL8 ( .A(N_13), .B(N_12), .C(GND), .D(GND), .Q(N_17), .S(N_11), .T(N_22) );
buff QL9 ( .A(N_8), .Q(N_24) );
xor2p QL10 ( .A(N_24), .B(N_25), .Q(Q[2]) );
xor2p QL11 ( .A(N_19), .B(N_23), .Q(Q[4]) );
mux2x2 QL12 ( .A(N_1), .B(N_1), .Q(N_15), .S(N_2) );
mux2x1 QL13 ( .A(N_1), .B(N_1), .Q(N_16), .S(N_3) );
and2i1 QL14 ( .A(A[0]), .B(B[0]), .Q(N_9) );
csblow QL15 ( .A0(A[0]), .A1(A[1]), .A1T(N_7), .B0(B[0]), .B1(B[1]), .C0_n(N_28),
           .C1(N_8) );
csbbitb QL16 ( .A(A[2]), .B(B[2]), .C0(N_5), .C1(N_6), .S0(N_25) );
csbbitb QL17 ( .A(A[3]), .B(B[3]), .C0(N_26), .C1(N_27), .S0(N_4) );
csbbita QL18 ( .A(A[4]), .B(B[4]), .C0(N_10), .C1(N_11), .S0(N_23) );
csbbita QL19 ( .A(A[5]), .B(B[5]), .C0(N_13), .C1(N_12), .S0(N_14) );
csbbita QL20 ( .A(A[6]), .B(B[6]), .C0(N_2), .C1(N_3), .S0(N_18) );
csbbita QL21 ( .A(A[7]), .B(B[7]), .S0(N_1) );
nand2i2 QL22 ( .A(N_28), .B(N_9), .Q(Q[0]) );

endmodule // sub8

`endif

`ifdef sub4
`else
`define sub4
module sub4( A , B, Q );
 input [3:0] A;
 input [3:0] B;
 output [3:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;

csamuxd QL1 ( .A(N_1), .Q(Q[3]), .S00(N_2), .S01(N_3), .S1(N_5) );
mux4x6 QL2 ( .A(N_8), .B(N_8), .C(N_8), .D(N_8), .Q(Q[1]), .S0(N_4), .S1(B[1]) );
xor2p QL3 ( .A(N_5), .B(N_7), .Q(Q[2]) );
and2i1 QL4 ( .A(A[0]), .B(B[0]), .Q(N_6) );
csblow QL5 ( .A0(A[0]), .A1(A[1]), .A1T(N_4), .B0(B[0]), .B1(B[1]), .C0_n(N_8),
          .C1(N_5) );
csbbitb QL6 ( .A(A[2]), .B(B[2]), .C0(N_2), .C1(N_3), .S0(N_7) );
csbbitb QL7 ( .A(A[3]), .B(B[3]), .S0(N_1) );
nand2i2 QL8 ( .A(N_8), .B(N_6), .Q(Q[0]) );

endmodule // sub4

`endif

`ifdef sub32
`else
`define sub32
module sub32( A , B, Q );
 input [31:0] A;
 input [31:0] B;
 output [31:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;
wire N_15;
wire N_16;
wire N_17;
wire N_18;
wire N_19;
wire N_20;
wire N_21;
wire N_22;
wire N_23;
wire N_24;
wire N_25;
wire N_26;
wire N_27;
wire N_28;
wire N_29;
wire N_30;
wire N_31;
wire N_32;
wire N_33;
wire N_34;
wire N_35;
wire N_36;
wire N_37;
wire N_38;
wire N_39;
wire N_40;
wire N_41;
wire N_42;
wire N_43;
wire N_44;
wire N_45;
wire N_46;
wire N_47;
wire N_48;
wire N_49;
wire N_50;
wire N_51;
wire N_52;
wire N_53;
wire N_54;
wire N_55;
wire N_56;
wire N_57;
wire N_58;
wire N_59;
wire N_60;
wire N_61;
wire N_62;
wire N_63;
wire N_64;
wire N_65;
wire N_66;
wire N_67;
wire N_68;
wire N_69;
wire N_70;
wire N_71;
wire N_72;
wire N_73;
wire N_74;
wire N_75;
wire N_76;
wire N_77;
wire N_78;
wire N_79;
wire N_80;
wire N_81;
wire N_82;
wire N_83;
wire N_84;
wire N_85;
wire N_86;
wire N_87;
wire N_88;
wire N_89;
wire N_90;
wire N_91;
wire N_92;
wire N_93;
wire N_94;
wire N_95;
wire N_96;
wire N_97;
wire N_98;
wire N_99;
wire N_100;
wire N_101;
wire N_102;
wire N_103;
wire N_104;
wire N_105;
wire N_106;
wire N_107;
wire N_108;
wire N_109;
wire N_110;
wire N_111;
wire N_112;
wire N_113;
wire N_114;
wire N_115;
wire N_116;
wire N_117;
wire N_118;
wire N_119;
wire N_120;
wire N_121;
wire N_122;
wire N_123;
wire N_124;
wire N_125;
wire N_126;
wire N_127;
wire N_128;
wire N_129;
wire N_130;
wire N_131;
wire N_132;
wire N_133;
wire N_134;
wire N_135;
wire N_136;
wire N_137;
wire N_138;
wire N_139;
wire N_140;
wire N_141;
wire N_142;
wire N_143;
wire N_144;
wire N_145;
wire N_146;
wire N_147;
wire N_148;
wire N_149;
wire N_150;
wire N_151;
wire N_152;
wire N_153;
wire N_154;
wire N_155;
wire N_156;
wire N_157;
wire N_158;
wire N_159;
wire N_160;
wire N_161;
wire N_162;
wire N_163;
wire N_164;
wire N_165;
wire N_166;
wire N_167;
wire N_168;
wire N_169;
wire N_170;
wire N_171;
wire N_172;
wire N_173;
wire N_174;
wire N_175;
wire N_176;
wire N_177;
wire N_178;
wire N_179;
wire N_180;
wire N_181;
wire N_182;
wire N_183;
wire N_184;
wire N_185;
wire N_186;
wire N_187;
wire N_188;
wire N_189;
wire C15A;
wire C15B;
wire N_190;
wire N_191;
wire N_192;
wire N_193;
wire N_194;
wire N_195;
wire N_196;
wire N_197;
wire C15C;
wire C15D;
wire N_198;
wire N_199;
wire N_200;
wire N_201;

mux2dxy QL1 ( .A(N_52), .B(N_52), .C(N_53), .D(N_53), .Q(N_50), .R(N_49), .S(N_51) );
xnor2p QL2 ( .A(A[31]), .B(B[31]), .Q(N_51) );
xor2p QL3 ( .A(C15A), .B(N_73), .Q(Q[16]) );
xor2p QL4 ( .A(N_138), .B(N_145), .Q(Q[8]) );
xor2p QL5 ( .A(N_111), .B(N_116), .Q(Q[4]) );
xor2p QL6 ( .A(N_115), .B(N_114), .Q(Q[2]) );
buff QL7 ( .A(N_120), .Q(N_111) );
buff QL8 ( .A(N_133), .Q(N_115) );
muxc2dx2 QL9 ( .A(N_128), .B(N_129), .C(N_128), .D(N_129), .Q(N_188), .R(N_124),
            .S(N_130), .T(N_117) );
muxb2dx2 QL10 ( .A(N_128), .B(N_129), .C(N_128), .D(N_129), .Q(N_189), .R(N_118),
             .S(N_131), .T(N_119) );
mux4x6 QL11 ( .A(N_201), .B(N_201), .C(N_201), .D(N_201), .Q(Q[1]), .S0(N_134),
           .S1(B[1]) );
csamuxd QL12 ( .A(N_127), .Q(Q[5]), .S00(N_119), .S01(N_117), .S1(N_111) );
csamuxd QL13 ( .A(N_137), .Q(Q[3]), .S00(N_136), .S01(N_135), .S1(N_115) );
csamuxc QL14 ( .A(N_113), .B(N_112), .Q(N_120), .S00(N_136), .S01(N_135),
            .S1(N_133) );
csamuxb QL15 ( .A(N_93), .B(N_81), .Q(Q[23]), .S00(N_77), .S01(N_78), .S1(C15B) );
csamuxb QL16 ( .A(N_94), .B(N_80), .Q(Q[22]), .S00(N_77), .S01(N_78), .S1(C15B) );
csamuxb QL17 ( .A(N_95), .B(N_96), .Q(Q[21]), .S00(N_77), .S01(N_78), .S1(C15B) );
csamuxb QL18 ( .A(N_55), .B(N_56), .Q(Q[25]), .S00(N_99), .S01(N_88), .S1(C15C) );
csamuxb QL19 ( .A(N_72), .B(N_71), .Q(Q[26]), .S00(N_99), .S01(N_88), .S1(C15C) );
csamuxb QL20 ( .A(N_58), .B(N_62), .Q(Q[27]), .S00(N_99), .S01(N_88), .S1(C15C) );
csamuxb QL21 ( .A(N_101), .B(N_103), .Q(Q[28]), .S00(N_110), .S01(N_109),
            .S1(C15D) );
csamuxb QL22 ( .A(N_102), .B(N_104), .Q(Q[29]), .S00(N_110), .S01(N_109),
            .S1(C15D) );
csamuxb QL23 ( .A(N_105), .B(N_107), .Q(Q[30]), .S00(N_110), .S01(N_109),
            .S1(C15D) );
csamuxb QL24 ( .A(N_106), .B(N_108), .Q(Q[31]), .S00(N_110), .S01(N_109),
            .S1(C15D) );
csamuxb QL25 ( .A(N_86), .B(N_84), .Q(Q[19]), .S00(N_83), .S01(N_82), .S1(C15A) );
csamuxb QL26 ( .A(N_100), .B(N_98), .Q(N_88), .S00(N_1), .S01(N_87), .S1(N_3) );
csamuxb QL27 ( .A(N_100), .B(N_98), .Q(N_99), .S00(N_1), .S01(N_87), .S1(N_2) );
csamuxb QL28 ( .A(N_100), .B(N_98), .Q(N_110), .S00(N_1), .S01(N_87), .S1(N_2) );
csamuxb QL29 ( .A(N_100), .B(N_98), .Q(N_109), .S00(N_1), .S01(N_87), .S1(N_3) );
csamuxb QL30 ( .A(N_123), .B(N_122), .Q(N_139), .S00(N_118), .S01(N_124),
            .S1(N_120) );
csamuxb QL31 ( .A(N_123), .B(N_122), .Q(N_138), .S00(N_189), .S01(N_188),
            .S1(N_120) );
csamuxb QL32 ( .A(N_192), .B(N_193), .Q(Q[13]), .S00(N_183), .S01(N_187),
            .S1(N_138) );
csamuxb QL33 ( .A(N_126), .B(N_125), .Q(Q[7]), .S00(N_189), .S01(N_188),
            .S1(N_111) );
csamuxb QL34 ( .A(N_197), .B(N_180), .Q(C15A), .S00(N_184), .S01(N_186),
            .S1(N_139) );
csamuxb QL35 ( .A(N_196), .B(N_181), .Q(Q[15]), .S00(N_183), .S01(N_187),
            .S1(N_138) );
csamuxb QL36 ( .A(N_194), .B(N_195), .Q(Q[14]), .S00(N_183), .S01(N_187),
            .S1(N_138) );
csamuxb QL37 ( .A(N_179), .B(N_178), .Q(Q[11]), .S00(N_182), .S01(N_190),
            .S1(N_138) );
csamuxb QL38 ( .A(N_197), .B(N_180), .Q(C15B), .S00(N_184), .S01(N_186),
            .S1(N_139) );
csamuxb QL39 ( .A(N_199), .B(N_200), .Q(C15C), .S00(N_184), .S01(N_186),
            .S1(N_139) );
csamuxb QL40 ( .A(N_199), .B(N_200), .Q(C15D), .S00(N_184), .S01(N_186),
            .S1(N_139) );
csamuxa QL41 ( .A(N_85), .Q(Q[18]), .S00(N_83), .S01(N_82), .S1(C15A) );
csamuxa QL42 ( .A(N_97), .Q(Q[20]), .S00(N_77), .S01(N_78), .S1(C15B) );
csamuxa QL43 ( .A(N_89), .Q(Q[24]), .S00(N_99), .S01(N_88), .S1(C15C) );
csamuxa QL44 ( .A(N_174), .Q(Q[10]), .S00(N_182), .S01(N_190), .S1(N_138) );
csamuxa QL45 ( .A(N_121), .Q(Q[6]), .S00(N_189), .S01(N_188), .S1(N_111) );
csamuxa QL46 ( .A(N_191), .Q(Q[12]), .S00(N_183), .S01(N_187), .S1(N_138) );
muxb2dx0 QL47 ( .A(N_74), .B(N_75), .C(N_74), .D(N_75), .Q(N_77), .R(N_2), .S(N_4),
             .T(N_83) );
muxb2dx0 QL48 ( .A(N_74), .B(N_75), .C(N_74), .D(N_75), .Q(N_78), .R(N_3), .S(N_76),
             .T(N_82) );
muxb2dx0 QL49 ( .A(N_15), .B(N_17), .C(N_18), .D(N_19), .Q(N_58), .R(N_59),
             .S(N_16), .T(N_57) );
muxb2dx0 QL50 ( .A(N_15), .B(N_17), .C(N_18), .D(N_19), .Q(N_62), .R(N_63),
             .S(N_20), .T(N_61) );
muxb2dx0 QL51 ( .A(N_175), .B(N_185), .C(N_175), .D(N_185), .Q(N_183), .R(N_184),
             .S(N_176), .T(N_182) );
muxb2dx0 QL52 ( .A(N_175), .B(N_185), .C(N_175), .D(N_185), .Q(N_187), .R(N_186),
             .S(N_177), .T(N_190) );
mux2x0 QL53 ( .A(N_54), .B(N_79), .Q(Q[17]), .S(C15A) );
mux2x0 QL54 ( .A(N_146), .B(N_147), .Q(Q[9]), .S(N_138) );
mux2dxx QL55 ( .A(N_92), .B(N_92), .C(N_90), .D(N_91), .Q(N_80), .R(N_81), .S(N_87) );
mux2dxx QL56 ( .A(N_48), .B(N_48), .C(N_50), .D(N_49), .Q(N_67), .R(N_68), .S(N_31) );
mux2dxx QL57 ( .A(N_48), .B(N_48), .C(N_50), .D(N_49), .Q(N_69), .R(N_70), .S(N_32) );
mux2dxx QL58 ( .A(N_64), .B(N_64), .C(N_65), .D(N_66), .Q(N_101), .R(N_102),
            .S(N_59) );
mux2dxx QL59 ( .A(N_64), .B(N_64), .C(N_65), .D(N_66), .Q(N_103), .R(N_104),
            .S(N_63) );
mux2dxx QL60 ( .A(N_92), .B(N_92), .C(N_90), .D(N_91), .Q(N_94), .R(N_93), .S(N_1) );
mux2dxx QL61 ( .A(N_198), .B(N_198), .C(N_159), .D(N_158), .Q(N_195), .R(N_181),
            .S(N_163) );
mux2dxx QL62 ( .A(N_198), .B(N_198), .C(N_159), .D(N_158), .Q(N_194), .R(N_196),
            .S(N_162) );
muxi2dx2 QL63 ( .A(N_5), .B(N_5), .C(N_7), .D(N_9), .Q(N_84), .R(N_75), .S(N_13) );
muxi2dx2 QL64 ( .A(N_6), .B(N_6), .C(N_8), .D(N_11), .Q(N_79), .R(N_76), .S(N_14) );
muxi2dx2 QL65 ( .A(N_21), .B(N_21), .C(N_23), .D(N_25), .Q(N_17), .R(N_19),
             .S(N_29) );
muxi2dx2 QL66 ( .A(N_22), .B(N_22), .C(N_24), .D(N_27), .Q(N_56), .R(N_20),
             .S(N_30) );
muxi2dx2 QL67 ( .A(N_33), .B(N_33), .C(N_34), .D(N_35), .Q(N_66), .R(N_32),
             .S(N_37) );
muxi2dx2 QL68 ( .A(N_38), .B(N_38), .C(N_40), .D(N_42), .Q(N_91), .R(N_98),
             .S(N_46) );
muxi2dx2 QL69 ( .A(N_39), .B(N_39), .C(N_41), .D(N_44), .Q(N_96), .R(N_87),
             .S(N_47) );
muxi2dx2 QL70 ( .A(N_144), .B(N_144), .C(N_143), .D(N_142), .Q(N_125), .R(N_122),
             .S(N_140) );
muxi2dx2 QL71 ( .A(N_148), .B(N_148), .C(N_150), .D(N_152), .Q(N_178), .R(N_185),
             .S(N_156) );
muxi2dx2 QL72 ( .A(N_149), .B(N_149), .C(N_151), .D(N_154), .Q(N_147), .R(N_177),
             .S(N_157) );
muxi2dx2 QL73 ( .A(N_164), .B(N_164), .C(N_166), .D(N_168), .Q(N_158), .R(N_160),
             .S(N_172) );
muxi2dx2 QL74 ( .A(N_165), .B(N_165), .C(N_167), .D(N_170), .Q(N_193), .R(N_163),
             .S(N_173) );
mux2dx2 QL75 ( .A(N_5), .B(N_5), .C(N_7), .D(N_9), .Q(N_86), .R(N_74), .S(N_10) );
mux2dx2 QL76 ( .A(N_6), .B(N_6), .C(N_8), .D(N_11), .Q(N_54), .R(N_4), .S(N_12) );
mux2dx2 QL77 ( .A(N_21), .B(N_21), .C(N_23), .D(N_25), .Q(N_15), .R(N_18), .S(N_26) );
mux2dx2 QL78 ( .A(N_22), .B(N_22), .C(N_24), .D(N_27), .Q(N_55), .R(N_16), .S(N_28) );
mux2dx2 QL79 ( .A(N_33), .B(N_33), .C(N_34), .D(N_35), .Q(N_65), .R(N_31), .S(N_36) );
mux2dx2 QL80 ( .A(N_38), .B(N_38), .C(N_40), .D(N_42), .Q(N_90), .R(N_100),
            .S(N_43) );
mux2dx2 QL81 ( .A(N_39), .B(N_39), .C(N_41), .D(N_44), .Q(N_95), .R(N_1), .S(N_45) );
mux2dx2 QL82 ( .A(N_57), .B(N_57), .C(N_61), .D(N_61), .Q(N_72), .R(N_71), .S(N_60) );
mux2dx2 QL83 ( .A(N_144), .B(N_144), .C(N_143), .D(N_142), .Q(N_126), .R(N_123),
            .S(N_141) );
mux2dx2 QL84 ( .A(N_148), .B(N_148), .C(N_150), .D(N_152), .Q(N_179), .R(N_175),
            .S(N_153) );
mux2dx2 QL85 ( .A(N_149), .B(N_149), .C(N_151), .D(N_154), .Q(N_146), .R(N_176),
            .S(N_155) );
mux2dx2 QL86 ( .A(N_164), .B(N_164), .C(N_166), .D(N_168), .Q(N_159), .R(N_161),
            .S(N_169) );
mux2dx2 QL87 ( .A(N_165), .B(N_165), .C(N_167), .D(N_170), .Q(N_192), .R(N_162),
            .S(N_171) );
mux2dx0 QL88 ( .A(N_67), .B(N_69), .C(N_68), .D(N_70), .Q(N_105), .R(N_106),
            .S(N_59) );
mux2dx0 QL89 ( .A(N_67), .B(N_69), .C(N_68), .D(N_70), .Q(N_107), .R(N_108),
            .S(N_63) );
mux2dx0 QL90 ( .A(N_161), .B(N_160), .C(N_161), .D(N_160), .Q(N_197), .R(N_199),
            .S(N_162) );
mux2dx0 QL91 ( .A(N_161), .B(N_160), .C(N_161), .D(N_160), .Q(N_180), .R(N_200),
            .S(N_163) );
csblow QL92 ( .A0(A[0]), .A1(A[1]), .A1T(N_134), .B0(B[0]), .B1(B[1]),
           .C0_n(N_201), .C1(N_133) );
and2i1 QL93 ( .A(A[0]), .B(B[0]), .Q(N_132) );
csbbitb QL94 ( .A(A[2]), .B(B[2]), .C0(N_136), .C1(N_135), .S0(N_114) );
csbbitb QL95 ( .A(A[3]), .B(B[3]), .C0(N_113), .C1(N_112), .S0(N_137) );
csbbita QL96 ( .A(A[16]), .B(B[16]), .C0(N_12), .C1(N_14), .S0(N_73) );
csbbita QL97 ( .A(A[17]), .B(B[17]), .C0(N_8), .C1(N_11), .S0(N_6) );
csbbita QL98 ( .A(A[18]), .B(B[18]), .C0(N_10), .C1(N_13), .S0(N_85) );
csbbita QL99 ( .A(A[19]), .B(B[19]), .C0(N_7), .C1(N_9), .S0(N_5) );
csbbita QL101 ( .A(A[20]), .B(B[20]), .C0(N_45), .C1(N_47), .S0(N_97) );
csbbita QL102 ( .A(A[21]), .B(B[21]), .C0(N_41), .C1(N_44), .S0(N_39) );
csbbita QL103 ( .A(A[22]), .B(B[22]), .C0(N_43), .C1(N_46), .S0(N_92) );
csbbita QL104 ( .A(A[23]), .B(B[23]), .C0(N_40), .C1(N_42), .S0(N_38) );
csbbita QL105 ( .A(A[24]), .B(B[24]), .C0(N_28), .C1(N_30), .S0(N_89) );
csbbita QL106 ( .A(A[25]), .B(B[25]), .C0(N_24), .C1(N_27), .S0(N_22) );
csbbita QL107 ( .A(A[26]), .B(B[26]), .C0(N_26), .C1(N_29), .S0(N_60) );
csbbita QL108 ( .A(A[27]), .B(B[27]), .C0(N_23), .C1(N_25), .S0(N_21) );
csbbita QL109 ( .A(A[28]), .B(B[28]), .C0(N_36), .C1(N_37), .S0(N_64) );
csbbita QL110 ( .A(A[29]), .B(B[29]), .C0(N_34), .C1(N_35), .S0(N_33) );
csbbita QL111 ( .A(A[30]), .B(B[30]), .C0(N_52), .C1(N_53), .S0(N_48) );
csbbita QL112 ( .A(A[4]), .B(B[4]), .C0(N_131), .C1(N_130), .S0(N_116) );
csbbita QL113 ( .A(A[5]), .B(B[5]), .C0(N_128), .C1(N_129), .S0(N_127) );
csbbita QL114 ( .A(A[6]), .B(B[6]), .C0(N_141), .C1(N_140), .S0(N_121) );
csbbita QL115 ( .A(A[7]), .B(B[7]), .C0(N_143), .C1(N_142), .S0(N_144) );
csbbita QL116 ( .A(A[8]), .B(B[8]), .C0(N_155), .C1(N_157), .S0(N_145) );
csbbita QL117 ( .A(A[9]), .B(B[9]), .C0(N_151), .C1(N_154), .S0(N_149) );
csbbita QL118 ( .A(A[10]), .B(B[10]), .C0(N_153), .C1(N_156), .S0(N_174) );
csbbita QL119 ( .A(A[11]), .B(B[11]), .C0(N_150), .C1(N_152), .S0(N_148) );
csbbita QL120 ( .A(A[12]), .B(B[12]), .C0(N_171), .C1(N_173), .S0(N_191) );
csbbita QL121 ( .A(A[13]), .B(B[13]), .C0(N_167), .C1(N_170), .S0(N_165) );
csbbita QL122 ( .A(A[14]), .B(B[14]), .C0(N_169), .C1(N_172), .S0(N_198) );
csbbita QL123 ( .A(A[15]), .B(B[15]), .C0(N_166), .C1(N_168), .S0(N_164) );
nand2i2 QL124 ( .A(N_201), .B(N_132), .Q(Q[0]) );

endmodule // sub32

`endif

`ifdef sub16
`else
`define sub16
module sub16( A , B, Q );
 input [15:0] A;
 input [15:0] B;
 output [15:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;
wire N_15;
wire N_16;
wire N_17;
wire N_18;
wire N_19;
wire N_20;
wire N_21;
wire N_22;
wire N_23;
wire N_24;
wire N_25;
wire N_26;
wire N_27;
wire N_28;
wire N_29;
wire N_30;
wire N_31;
wire N_32;
wire N_33;
wire N_34;
wire N_35;
wire N_36;
wire N_37;
wire N_38;
wire N_39;
wire N_40;
wire N_41;
wire N_42;
wire N_43;
wire N_44;
wire N_45;
wire N_46;
wire N_47;
wire N_48;
wire N_49;
wire N_50;
wire N_51;
wire N_52;
wire N_53;
wire N_54;
wire N_55;
wire N_56;
wire N_57;
wire N_58;
wire N_59;
wire N_60;
wire N_61;
wire N_62;
wire N_63;
wire N_64;
wire N_65;
wire N_66;
wire N_67;
wire N_68;
wire N_69;
wire N_70;
wire N_71;
wire N_72;
wire N_73;
wire N_74;
wire N_75;
wire N_76;
wire N_77;
wire N_78;
wire N_79;
wire N_80;
wire N_81;
wire N_82;
wire N_83;

mux2dx2 QL1 ( .A(N_12), .B(N_12), .C(N_16), .D(N_23), .Q(N_60), .R(N_65), .S(N_24) );
mux2dx2 QL2 ( .A(N_11), .B(N_11), .C(N_15), .D(N_21), .Q(N_33), .R(N_4), .S(N_22) );
mux2dx2 QL3 ( .A(N_10), .B(N_10), .C(N_14), .D(N_19), .Q(N_3), .R(N_6), .S(N_20) );
mux2dx2 QL4 ( .A(N_9), .B(N_9), .C(N_13), .D(N_17), .Q(N_43), .R(N_2), .S(N_18) );
muxi2dx2 QL5 ( .A(N_12), .B(N_12), .C(N_16), .D(N_23), .Q(N_61), .R(N_66), .S(N_28) );
muxi2dx2 QL6 ( .A(N_11), .B(N_11), .C(N_15), .D(N_21), .Q(N_34), .R(N_8), .S(N_27) );
muxi2dx2 QL7 ( .A(N_10), .B(N_10), .C(N_14), .D(N_19), .Q(N_5), .R(N_7), .S(N_26) );
muxi2dx2 QL8 ( .A(N_9), .B(N_9), .C(N_13), .D(N_17), .Q(N_44), .R(N_29), .S(N_25) );
mux2dxx QL9 ( .A(N_1), .B(N_1), .C(N_79), .D(N_78), .Q(N_45), .R(N_46), .S(N_2) );
mux2dxx QL10 ( .A(N_1), .B(N_1), .C(N_79), .D(N_78), .Q(N_47), .R(N_48), .S(N_29) );
mux2x0 QL11 ( .A(N_33), .B(N_34), .Q(Q[9]), .S(N_31) );
mux2x0 QL12 ( .A(N_36), .B(N_40), .Q(Q[11]), .S(N_31) );
muxb2dx0 QL13 ( .A(N_3), .B(N_5), .C(N_6), .D(N_7), .Q(N_36), .R(N_37), .S(N_4),
             .T(N_35) );
muxb2dx0 QL14 ( .A(N_3), .B(N_5), .C(N_6), .D(N_7), .Q(N_40), .R(N_41), .S(N_8),
             .T(N_39) );
csamuxa QL15 ( .A(N_67), .Q(Q[6]), .S00(N_70), .S01(N_63), .S1(N_82) );
csamuxa QL16 ( .A(N_42), .Q(Q[12]), .S00(N_37), .S01(N_41), .S1(N_30) );
csamuxa QL17 ( .A(N_38), .Q(Q[10]), .S00(N_35), .S01(N_39), .S1(N_31) );
csamuxb QL18 ( .A(N_60), .B(N_61), .Q(Q[7]), .S00(N_70), .S01(N_63), .S1(N_82) );
csamuxb QL19 ( .A(N_43), .B(N_44), .Q(Q[13]), .S00(N_37), .S01(N_41), .S1(N_30) );
csamuxb QL20 ( .A(N_45), .B(N_47), .Q(Q[14]), .S00(N_37), .S01(N_41), .S1(N_30) );
csamuxb QL21 ( .A(N_46), .B(N_48), .Q(Q[15]), .S00(N_37), .S01(N_41), .S1(N_30) );
csamuxb QL22 ( .A(N_65), .B(N_66), .Q(N_31), .S00(N_62), .S01(N_64), .S1(N_68) );
csamuxb QL23 ( .A(N_65), .B(N_66), .Q(N_30), .S00(N_62), .S01(N_64), .S1(N_68) );
csamuxc QL24 ( .A(N_80), .B(N_81), .Q(N_68), .S00(N_50), .S01(N_51), .S1(N_53) );
csamuxd QL25 ( .A(N_49), .Q(Q[3]), .S00(N_50), .S01(N_51), .S1(N_73) );
csamuxd QL26 ( .A(N_59), .Q(Q[5]), .S00(N_69), .S01(N_71), .S1(N_82) );
mux4x6 QL27 ( .A(N_83), .B(N_83), .C(N_83), .D(N_83), .Q(Q[1]), .S0(N_52),
           .S1(B[1]) );
muxb2dx2 QL28 ( .A(N_58), .B(N_57), .C(N_58), .D(N_57), .Q(N_70), .R(N_62),
             .S(N_55), .T(N_69) );
muxc2dx2 QL29 ( .A(N_58), .B(N_57), .C(N_58), .D(N_57), .Q(N_63), .R(N_64),
             .S(N_56), .T(N_71) );
buff QL30 ( .A(N_53), .Q(N_73) );
buff QL31 ( .A(N_68), .Q(N_82) );
xor2p QL32 ( .A(N_73), .B(N_74), .Q(Q[2]) );
xor2p QL33 ( .A(N_82), .B(N_72), .Q(Q[4]) );
xor2p QL34 ( .A(N_31), .B(N_32), .Q(Q[8]) );
mux2dxy QL35 ( .A(N_75), .B(N_75), .C(N_76), .D(N_76), .Q(N_79), .R(N_78), .S(N_77) );
csblow QL36 ( .A0(A[0]), .A1(A[1]), .A1T(N_52), .B0(B[0]), .B1(B[1]), .C0_n(N_83),
           .C1(N_53) );
and2i1 QL37 ( .A(A[0]), .B(B[0]), .Q(N_54) );
csbbitb QL38 ( .A(A[2]), .B(B[2]), .C0(N_50), .C1(N_51), .S0(N_74) );
csbbitb QL39 ( .A(A[3]), .B(B[3]), .C0(N_80), .C1(N_81), .S0(N_49) );
csbbita QL40 ( .A(A[4]), .B(B[4]), .C0(N_55), .C1(N_56), .S0(N_72) );
csbbita QL41 ( .A(A[5]), .B(B[5]), .C0(N_58), .C1(N_57), .S0(N_59) );
csbbita QL42 ( .A(A[6]), .B(B[6]), .C0(N_24), .C1(N_28), .S0(N_67) );
csbbita QL43 ( .A(A[7]), .B(B[7]), .C0(N_16), .C1(N_23), .S0(N_12) );
csbbita QL44 ( .A(A[8]), .B(B[8]), .C0(N_22), .C1(N_27), .S0(N_32) );
csbbita QL45 ( .A(A[9]), .B(B[9]), .C0(N_15), .C1(N_21), .S0(N_11) );
csbbita QL46 ( .A(A[10]), .B(B[10]), .C0(N_20), .C1(N_26), .S0(N_38) );
csbbita QL47 ( .A(A[11]), .B(B[11]), .C0(N_14), .C1(N_19), .S0(N_10) );
csbbita QL48 ( .A(A[12]), .B(B[12]), .C0(N_18), .C1(N_25), .S0(N_42) );
csbbita QL49 ( .A(A[13]), .B(B[13]), .C0(N_13), .C1(N_17), .S0(N_9) );
csbbita QL50 ( .A(A[14]), .B(B[14]), .C0(N_75), .C1(N_76), .S0(N_1) );
xnor2p QL51 ( .A(A[15]), .B(B[15]), .Q(N_77) );
nand2i2 QL52 ( .A(N_83), .B(N_54), .Q(Q[0]) );

endmodule // sub16

`endif

`ifdef radd8
`else
`define radd8
module radd8( A , B, CI, CO, S );
 input [7:0] A;
 input [7:0] B;
input CI;
output CO;
 output [7:0] S;
wire N_1;

radd4 QL2 ( .A({ A[7:4] }), .B({ B[7:4] }), .CI(N_1), .CO(CO), .S({ S[7:4] }) );
radd4 QL1 ( .A({ A[3:0] }), .B({ B[3:0] }), .CI(CI), .CO(N_1), .S({ S[3:0] }) );

endmodule // radd8

`endif

`ifdef radd4
`else
`define radd4
module radd4( A , B, CI, CO, S );
 input [3:0] A;
 input [3:0] B;
input CI;
output CO;
 output [3:0] S;
wire N_1;
wire N_2;
wire N_3;

fadd1 QL1 ( .A(A[0]), .B(B[0]), .CI(CI), .CO(N_1), .S(S[0]) );
fadd1 QL2 ( .A(A[1]), .B(B[1]), .CI(N_1), .CO(N_2), .S(S[1]) );
fadd1 QL3 ( .A(A[2]), .B(B[2]), .CI(N_2), .CO(N_3), .S(S[2]) );
fadd1 QL4 ( .A(A[3]), .B(B[3]), .CI(N_3), .CO(CO), .S(S[3]) );

endmodule // radd4

`endif

`ifdef radd16
`else
`define radd16
module radd16( A , B, CI, CO, S );
 input [15:0] A;
 input [15:0] B;
input CI;
output CO;
 output [15:0] S;
wire N_1;
wire N_2;
wire N_3;

radd4 QL4 ( .A({ A[15:12] }), .B({ B[15:12] }), .CI(N_1), .CO(CO),
         .S({ S[15:12] }) );
radd4 QL3 ( .A({ A[11:8] }), .B({ B[11:8] }), .CI(N_2), .CO(N_1), .S({ S[11:8] }) );
radd4 QL2 ( .A({ A[7:4] }), .B({ B[7:4] }), .CI(N_3), .CO(N_2), .S({ S[7:4] }) );
radd4 QL1 ( .A({ A[3:0] }), .B({ B[3:0] }), .CI(CI), .CO(N_3), .S({ S[3:0] }) );

endmodule // radd16

`endif

`ifdef mult4x4
`else
`define mult4x4
module mult4x4( X , Y, P );
 output [7:0] P;
 input [3:0] X;
 input [3:0] Y;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;
wire N_15;
wire N_16;
supply0 GND;

mbitc QL1 ( .A(N_7), .B0(Y[0]), .B1(X[2]), .CI(N_10), .CO(N_9), .S(P[2]) );
mbitc QL2 ( .A(N_8), .B0(Y[1]), .B1(X[2]), .CI(N_13), .CO(N_12), .S(N_5) );
mbitc QL3 ( .A(N_6), .B0(Y[1]), .B1(X[3]), .CI(N_12), .CO(N_11), .S(N_3) );
mbitc QL4 ( .A(N_5), .B0(Y[0]), .B1(X[3]), .CI(N_9), .CO(N_1), .S(P[3]) );
mbitc QL5 ( .A(N_4), .B0(N_3), .B1(N_1), .CI(N_11), .CO(N_2), .S(P[5]) );
mbitb QL6 ( .A0(Y[3]), .A1(X[3]), .B(N_2), .CI(N_14), .CO(P[7]), .S(P[6]) );
mbita QL7 ( .A0(Y[1]), .A1(X[0]), .B0(Y[0]), .B1(X[1]), .CI(GND), .CO(N_10),
         .S(P[1]) );
mbita QL8 ( .A0(Y[2]), .A1(X[0]), .B0(Y[1]), .B1(X[1]), .CI(GND), .CO(N_13),
         .S(N_7) );
mbita QL9 ( .A0(Y[3]), .A1(X[0]), .B0(Y[2]), .B1(X[1]), .CI(GND), .CO(N_16),
         .S(N_8) );
mbita QL10 ( .A0(Y[3]), .A1(X[1]), .B0(Y[2]), .B1(X[2]), .CI(N_16), .CO(N_15),
          .S(N_6) );
mbita QL11 ( .A0(Y[3]), .A1(X[2]), .B0(Y[2]), .B1(X[3]), .CI(N_15), .CO(N_14),
          .S(N_4) );
xor2i0 QL12 ( .A(N_3), .B(N_1), .Q(P[4]) );
and2i0 QL13 ( .A(Y[0]), .B(X[0]), .Q(P[0]) );

endmodule // mult4x4

`endif

`ifdef hadd1
`else
`define hadd1
module hadd1( A , B, CO, S );
input A, B;
output CO, S;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
supply1 VCC;

frag_m I_2 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(B), .D2(GND), .E1(VCC),
          .E2(B), .NS(N_1), .NZ(S), .OS(CO) );
frag_f I_1 ( .F1(A), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_a QL3 ( .A1(A), .A2(GND), .A3(B), .A4(GND), .A5(VCC), .A6(GND), .AZ(CO) );

endmodule // hadd1

`endif

`ifdef fadd1
`else
`define fadd1
module fadd1( A , B, CI, CO, S );
input A, B, CI;
output CO, S;

maj3i0 QL2 ( .A(A), .B(B), .C(CI), .Q(CO) );
xor3i0 QL1 ( .A(CI), .B(B), .C(A), .Q(S) );

endmodule // fadd1

`endif

`ifdef comp8
`else
`define comp8
module comp8( A , B, EQ );
 input [7:0] A;
 input [7:0] B;
output EQ;
parameter syn_macro = 1, ql_pack = 1;
wire N_1;
wire N_2;
supply0 GND;
supply1 VCC;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;

eqcombit QL1 ( .A1(A[0]), .A2(A[1]), .B1(B[0]), .B2(B[1]), .EQ1(N_4), .EQ2(N_2) );
eqcombit QL2 ( .A1(A[2]), .A2(A[3]), .B1(B[2]), .B2(B[3]), .EQ1(N_5), .EQ2(N_1) );
eqcombit QL3 ( .A1(A[4]), .A2(A[5]), .B1(B[4]), .B2(B[5]), .EQ1(N_6), .EQ2(N_3) );
eqcombit QL4 ( .A1(A[6]), .A2(A[7]), .B1(B[6]), .B2(B[7]), .EQ1(N_7), .EQ2(N_8) );
and14i7 QL5 ( .A(N_2), .B(N_1), .C(N_3), .D(N_8), .E(VCC), .F(VCC), .G(VCC), .H(GND),
           .I(N_4), .J(N_5), .K(N_6), .L(N_7), .M(GND), .N(GND), .Q(EQ) );

endmodule // comp8

`endif

`ifdef comp4
`else
`define comp4
module comp4( A , B, EQ );
 input [3:0] A;
 input [3:0] B;
output EQ;
parameter syn_macro = 1, ql_pack = 1;
wire N_1;
wire N_2;
wire N_3;
wire N_4;

eqcombit QL1 ( .A1(A[0]), .A2(A[1]), .B1(B[0]), .B2(B[1]), .EQ1(N_3), .EQ2(N_2) );
eqcombit QL2 ( .A1(A[2]), .A2(A[3]), .B1(B[2]), .B2(B[3]), .EQ1(N_4), .EQ2(N_1) );
and4i2 QL3 ( .A(N_2), .B(N_1), .C(N_3), .D(N_4), .Q(EQ) );

endmodule // comp4

`endif

`ifdef comp12
`else
`define comp12
module comp12( A , B, EQ );
 input [11:0] A;
 input [11:0] B;
output EQ;
parameter syn_macro = 1, ql_pack = 1;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
supply0 GND;
supply1 VCC;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;

eqcombit QL1 ( .A1(A[0]), .A2(A[1]), .B1(B[0]), .B2(B[1]), .EQ1(N_8), .EQ2(N_6) );
eqcombit QL2 ( .A1(A[2]), .A2(A[3]), .B1(B[2]), .B2(B[3]), .EQ1(N_9), .EQ2(N_5) );
eqcombit QL3 ( .A1(A[4]), .A2(A[5]), .B1(B[4]), .B2(B[5]), .EQ1(N_10), .EQ2(N_7) );
eqcombit QL4 ( .A1(A[6]), .A2(A[7]), .B1(B[6]), .B2(B[7]), .EQ1(N_11), .EQ2(N_12) );
eqcombit QL5 ( .A1(A[8]), .A2(A[9]), .B1(B[8]), .B2(B[9]), .EQ1(N_2), .EQ2(N_4) );
eqcombit QL6 ( .A1(A[10]), .A2(A[11]), .B1(B[10]), .B2(B[11]), .EQ1(N_1),
            .EQ2(N_3) );
and14i7 QL7 ( .A(N_6), .B(N_5), .C(N_7), .D(N_12), .E(N_4), .F(N_3), .G(VCC),
           .H(GND), .I(N_8), .J(N_9), .K(N_10), .L(N_11), .M(N_2), .N(N_1),
           .Q(EQ) );

endmodule // comp12

`endif

`ifdef add8
`else
`define add8
module add8( A , B, Q );
 input [7:0] A;
 input [7:0] B;
 output [7:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;
wire N_15;
wire N_16;
wire N_17;
wire N_18;
wire N_19;
wire N_20;
wire N_21;
wire N_22;
wire N_23;
wire N_24;
wire N_25;
wire N_26;
wire N_27;
wire N_28;
supply0 GND;

csamuxa QL1 ( .A(N_19), .Q(Q[6]), .S00(N_22), .S01(N_18), .S1(N_20) );
csamuxb QL2 ( .A(N_16), .B(N_17), .Q(Q[7]), .S00(N_22), .S01(N_18), .S1(N_20) );
csamuxc QL3 ( .A(N_27), .B(N_28), .Q(N_20), .S00(N_5), .S01(N_6), .S1(N_8) );
csamuxd QL4 ( .A(N_4), .Q(Q[3]), .S00(N_5), .S01(N_6), .S1(N_25) );
csamuxd QL5 ( .A(N_15), .Q(Q[5]), .S00(N_21), .S01(N_23), .S1(N_20) );
mux4x6 QL6 ( .A(N_10), .B(N_10), .C(N_10), .D(N_10), .Q(Q[1]), .S0(N_7), .S1(B[1]) );
csalow QL7 ( .A0(A[0]), .A1(A[1]), .A1T(N_7), .B0(B[0]), .B1(B[1]), .C0(N_10),
          .C1(N_8) );
and2i2 QL8 ( .A(N_9), .B(N_10), .Q(Q[0]) );
nor2i0 QL9 ( .A(B[0]), .B(A[0]), .Q(N_9) );
muxb2dx2 QL10 ( .A(N_14), .B(N_13), .C(GND), .D(GND), .Q(N_22), .S(N_11), .T(N_21) );
muxc2dx2 QL11 ( .A(N_14), .B(N_13), .C(GND), .D(GND), .Q(N_18), .S(N_12), .T(N_23) );
buff QL12 ( .A(N_8), .Q(N_25) );
csabita QL13 ( .A(A[4]), .B(B[4]), .C0(N_11), .C1(N_12), .S0(N_24) );
csabita QL14 ( .A(A[5]), .B(B[5]), .C0(N_14), .C1(N_13), .S0(N_15) );
csabita QL15 ( .A(A[6]), .B(B[6]), .C0(N_2), .C1(N_3), .S0(N_19) );
csabita QL16 ( .A(A[7]), .B(B[7]), .S0(N_1) );
csabitb QL17 ( .A(A[2]), .B(B[2]), .C0(N_5), .C1(N_6), .S0(N_26) );
csabitb QL18 ( .A(A[3]), .B(B[3]), .C0(N_27), .C1(N_28), .S0(N_4) );
xor2p QL19 ( .A(N_25), .B(N_26), .Q(Q[2]) );
xor2p QL20 ( .A(N_20), .B(N_24), .Q(Q[4]) );
mux2x2 QL21 ( .A(N_1), .B(N_1), .Q(N_16), .S(N_2) );
mux2x1 QL22 ( .A(N_1), .B(N_1), .Q(N_17), .S(N_3) );

endmodule // add8

`endif

`ifdef add4
`else
`define add4
module add4( A , B, Q );
 input [3:0] A;
 input [3:0] B;
 output [3:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;

csamuxd QL1 ( .A(N_1), .Q(Q[3]), .S00(N_2), .S01(N_3), .S1(N_5) );
mux4x6 QL2 ( .A(N_7), .B(N_7), .C(N_7), .D(N_7), .Q(Q[1]), .S0(N_4), .S1(B[1]) );
csalow QL3 ( .A0(A[0]), .A1(A[1]), .A1T(N_4), .B0(B[0]), .B1(B[1]), .C0(N_7),
          .C1(N_5) );
and2i2 QL4 ( .A(N_6), .B(N_7), .Q(Q[0]) );
nor2i0 QL5 ( .A(B[0]), .B(A[0]), .Q(N_6) );
csabitb QL6 ( .A(A[2]), .B(B[2]), .C0(N_2), .C1(N_3), .S0(N_8) );
csabitb QL7 ( .A(A[3]), .B(B[3]), .S0(N_1) );
xor2p QL8 ( .A(N_5), .B(N_8), .Q(Q[2]) );

endmodule // add4

`endif

`ifdef add32
`else
`define add32
module add32( A , B, Q );
 input [31:0] A;
 input [31:0] B;
 output [31:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;
wire N_15;
wire N_16;
wire N_17;
wire N_18;
wire N_19;
wire N_20;
wire N_21;
wire N_22;
wire N_23;
wire N_24;
wire N_25;
wire N_26;
wire N_27;
wire N_28;
wire N_29;
wire N_30;
wire N_31;
wire N_32;
wire N_33;
wire N_34;
wire N_35;
wire N_36;
wire N_37;
wire N_38;
wire N_39;
wire N_40;
wire N_41;
wire N_42;
wire N_43;
wire N_44;
wire N_45;
wire N_46;
wire N_47;
wire N_48;
wire N_49;
wire N_50;
wire N_51;
wire N_52;
wire N_53;
wire N_54;
wire N_55;
wire N_56;
wire N_57;
wire N_58;
wire N_59;
wire N_60;
wire N_61;
wire N_62;
wire N_63;
wire N_64;
wire N_65;
wire N_66;
wire N_67;
wire N_68;
wire N_69;
wire N_70;
wire N_71;
wire N_72;
wire N_73;
wire N_74;
wire N_75;
wire N_76;
wire N_77;
wire N_78;
wire N_79;
wire N_80;
wire N_81;
wire N_82;
wire N_83;
wire N_84;
wire N_85;
wire N_86;
wire N_87;
wire N_88;
wire N_89;
wire N_90;
wire N_91;
wire N_92;
wire N_93;
wire N_94;
wire N_95;
wire N_96;
wire N_97;
wire N_98;
wire N_99;
wire N_100;
wire N_101;
wire N_102;
wire N_103;
wire N_104;
wire N_105;
wire N_106;
wire N_107;
wire N_108;
wire N_109;
wire N_110;
wire N_111;
wire N_112;
wire N_113;
wire N_114;
wire N_115;
wire N_116;
wire N_117;
wire N_118;
wire N_119;
wire N_120;
wire N_121;
wire N_122;
wire N_123;
wire N_124;
wire N_125;
wire N_126;
wire N_127;
wire N_128;
wire N_129;
wire N_130;
wire N_131;
wire N_132;
wire N_133;
wire N_134;
wire N_135;
wire N_136;
wire N_137;
wire N_138;
wire N_139;
wire N_140;
wire N_141;
wire N_142;
wire N_143;
wire N_144;
wire N_145;
wire N_146;
wire N_147;
wire N_148;
wire N_149;
wire N_150;
wire N_151;
wire N_152;
wire N_153;
wire N_154;
wire N_155;
wire N_156;
wire N_157;
wire N_158;
wire N_159;
wire N_160;
wire N_161;
wire N_162;
wire N_163;
wire N_164;
wire N_165;
wire N_166;
wire N_167;
wire N_168;
wire N_169;
wire N_170;
wire N_171;
wire N_172;
wire N_173;
wire N_174;
wire N_175;
wire N_176;
wire N_177;
wire N_178;
wire N_179;
wire N_180;
wire N_181;
wire N_182;
wire N_183;
wire N_184;
wire N_185;
wire N_186;
wire N_187;
wire N_188;
wire N_189;
wire N_190;
wire C15A;
wire C15B;
wire N_191;
wire N_192;
wire N_193;
wire N_194;
wire N_195;
wire N_196;
wire N_197;
wire N_198;
wire C15C;
wire C15D;
wire N_199;
wire N_200;
wire N_201;

mux2dxy QL1 ( .A(N_52), .B(N_52), .C(N_53), .D(N_53), .Q(N_50), .R(N_49), .S(N_51) );
xor2p QL2 ( .A(A[31]), .B(B[31]), .Q(N_51) );
xor2p QL3 ( .A(C15A), .B(N_73), .Q(Q[16]) );
xor2p QL4 ( .A(N_139), .B(N_146), .Q(Q[8]) );
xor2p QL5 ( .A(N_111), .B(N_116), .Q(Q[4]) );
xor2p QL6 ( .A(N_115), .B(N_114), .Q(Q[2]) );
csabitb QL7 ( .A(A[3]), .B(B[3]), .C0(N_113), .C1(N_112), .S0(N_138) );
csabitb QL8 ( .A(A[2]), .B(B[2]), .C0(N_137), .C1(N_136), .S0(N_114) );
csabita QL9 ( .A(A[18]), .B(B[18]), .C0(N_10), .C1(N_13), .S0(N_85) );
csabita QL10 ( .A(A[19]), .B(B[19]), .C0(N_7), .C1(N_9), .S0(N_5) );
csabita QL11 ( .A(A[20]), .B(B[20]), .C0(N_45), .C1(N_47), .S0(N_97) );
csabita QL12 ( .A(A[21]), .B(B[21]), .C0(N_41), .C1(N_44), .S0(N_39) );
csabita QL13 ( .A(A[22]), .B(B[22]), .C0(N_43), .C1(N_46), .S0(N_92) );
csabita QL14 ( .A(A[23]), .B(B[23]), .C0(N_40), .C1(N_42), .S0(N_38) );
csabita QL15 ( .A(A[24]), .B(B[24]), .C0(N_28), .C1(N_30), .S0(N_89) );
csabita QL16 ( .A(A[25]), .B(B[25]), .C0(N_24), .C1(N_27), .S0(N_22) );
csabita QL17 ( .A(A[26]), .B(B[26]), .C0(N_26), .C1(N_29), .S0(N_60) );
csabita QL18 ( .A(A[27]), .B(B[27]), .C0(N_23), .C1(N_25), .S0(N_21) );
csabita QL19 ( .A(A[28]), .B(B[28]), .C0(N_36), .C1(N_37), .S0(N_64) );
csabita QL20 ( .A(A[29]), .B(B[29]), .C0(N_34), .C1(N_35), .S0(N_33) );
csabita QL21 ( .A(A[30]), .B(B[30]), .C0(N_52), .C1(N_53), .S0(N_48) );
csabita QL22 ( .A(A[17]), .B(B[17]), .C0(N_8), .C1(N_11), .S0(N_6) );
csabita QL23 ( .A(A[16]), .B(B[16]), .C0(N_12), .C1(N_14), .S0(N_73) );
csabita QL24 ( .A(A[14]), .B(B[14]), .C0(N_170), .C1(N_173), .S0(N_199) );
csabita QL25 ( .A(A[13]), .B(B[13]), .C0(N_168), .C1(N_171), .S0(N_166) );
csabita QL26 ( .A(A[12]), .B(B[12]), .C0(N_172), .C1(N_174), .S0(N_192) );
csabita QL27 ( .A(A[11]), .B(B[11]), .C0(N_151), .C1(N_153), .S0(N_149) );
csabita QL28 ( .A(A[10]), .B(B[10]), .C0(N_154), .C1(N_157), .S0(N_175) );
csabita QL29 ( .A(A[9]), .B(B[9]), .C0(N_152), .C1(N_155), .S0(N_150) );
csabita QL30 ( .A(A[8]), .B(B[8]), .C0(N_156), .C1(N_158), .S0(N_146) );
csabita QL31 ( .A(A[7]), .B(B[7]), .C0(N_144), .C1(N_143), .S0(N_145) );
csabita QL32 ( .A(A[6]), .B(B[6]), .C0(N_142), .C1(N_141), .S0(N_121) );
csabita QL33 ( .A(A[5]), .B(B[5]), .C0(N_128), .C1(N_129), .S0(N_127) );
csabita QL34 ( .A(A[4]), .B(B[4]), .C0(N_131), .C1(N_130), .S0(N_116) );
csabita QL35 ( .A(A[15]), .B(B[15]), .C0(N_167), .C1(N_169), .S0(N_165) );
buff QL36 ( .A(N_120), .Q(N_111) );
buff QL37 ( .A(N_134), .Q(N_115) );
muxc2dx2 QL38 ( .A(N_128), .B(N_129), .C(N_128), .D(N_129), .Q(N_189), .R(N_124),
             .S(N_130), .T(N_117) );
muxb2dx2 QL39 ( .A(N_128), .B(N_129), .C(N_128), .D(N_129), .Q(N_190), .R(N_118),
             .S(N_131), .T(N_119) );
nor2i0 QL40 ( .A(B[0]), .B(A[0]), .Q(N_133) );
and2i2 QL41 ( .A(N_133), .B(N_132), .Q(Q[0]) );
csalow QL42 ( .A0(A[0]), .A1(A[1]), .A1T(N_135), .B0(B[0]), .B1(B[1]), .C0(N_132),
           .C1(N_134) );
mux4x6 QL43 ( .A(N_132), .B(N_132), .C(N_132), .D(N_132), .Q(Q[1]), .S0(N_135),
           .S1(B[1]) );
csamuxd QL44 ( .A(N_127), .Q(Q[5]), .S00(N_119), .S01(N_117), .S1(N_111) );
csamuxd QL45 ( .A(N_138), .Q(Q[3]), .S00(N_137), .S01(N_136), .S1(N_115) );
csamuxc QL46 ( .A(N_113), .B(N_112), .Q(N_120), .S00(N_137), .S01(N_136),
            .S1(N_134) );
csamuxb QL47 ( .A(N_93), .B(N_81), .Q(Q[23]), .S00(N_77), .S01(N_78), .S1(C15B) );
csamuxb QL48 ( .A(N_94), .B(N_80), .Q(Q[22]), .S00(N_77), .S01(N_78), .S1(C15B) );
csamuxb QL49 ( .A(N_95), .B(N_96), .Q(Q[21]), .S00(N_77), .S01(N_78), .S1(C15B) );
csamuxb QL50 ( .A(N_55), .B(N_56), .Q(Q[25]), .S00(N_99), .S01(N_88), .S1(C15C) );
csamuxb QL51 ( .A(N_72), .B(N_71), .Q(Q[26]), .S00(N_99), .S01(N_88), .S1(C15C) );
csamuxb QL52 ( .A(N_58), .B(N_62), .Q(Q[27]), .S00(N_99), .S01(N_88), .S1(C15C) );
csamuxb QL53 ( .A(N_101), .B(N_103), .Q(Q[28]), .S00(N_110), .S01(N_109),
            .S1(C15D) );
csamuxb QL54 ( .A(N_102), .B(N_104), .Q(Q[29]), .S00(N_110), .S01(N_109),
            .S1(C15D) );
csamuxb QL55 ( .A(N_105), .B(N_107), .Q(Q[30]), .S00(N_110), .S01(N_109),
            .S1(C15D) );
csamuxb QL56 ( .A(N_106), .B(N_108), .Q(Q[31]), .S00(N_110), .S01(N_109),
            .S1(C15D) );
csamuxb QL57 ( .A(N_86), .B(N_84), .Q(Q[19]), .S00(N_83), .S01(N_82), .S1(C15A) );
csamuxb QL58 ( .A(N_100), .B(N_98), .Q(N_88), .S00(N_1), .S01(N_87), .S1(N_3) );
csamuxb QL59 ( .A(N_100), .B(N_98), .Q(N_99), .S00(N_1), .S01(N_87), .S1(N_2) );
csamuxb QL60 ( .A(N_100), .B(N_98), .Q(N_110), .S00(N_1), .S01(N_87), .S1(N_2) );
csamuxb QL61 ( .A(N_100), .B(N_98), .Q(N_109), .S00(N_1), .S01(N_87), .S1(N_3) );
csamuxb QL62 ( .A(N_123), .B(N_122), .Q(N_140), .S00(N_118), .S01(N_124),
            .S1(N_120) );
csamuxb QL63 ( .A(N_123), .B(N_122), .Q(N_139), .S00(N_190), .S01(N_189),
            .S1(N_120) );
csamuxb QL64 ( .A(N_193), .B(N_194), .Q(Q[13]), .S00(N_184), .S01(N_188),
            .S1(N_139) );
csamuxb QL65 ( .A(N_126), .B(N_125), .Q(Q[7]), .S00(N_190), .S01(N_189),
            .S1(N_111) );
csamuxb QL66 ( .A(N_198), .B(N_181), .Q(C15A), .S00(N_185), .S01(N_187),
            .S1(N_140) );
csamuxb QL67 ( .A(N_197), .B(N_182), .Q(Q[15]), .S00(N_184), .S01(N_188),
            .S1(N_139) );
csamuxb QL68 ( .A(N_195), .B(N_196), .Q(Q[14]), .S00(N_184), .S01(N_188),
            .S1(N_139) );
csamuxb QL69 ( .A(N_180), .B(N_179), .Q(Q[11]), .S00(N_183), .S01(N_191),
            .S1(N_139) );
csamuxb QL70 ( .A(N_198), .B(N_181), .Q(C15B), .S00(N_185), .S01(N_187),
            .S1(N_140) );
csamuxb QL71 ( .A(N_200), .B(N_201), .Q(C15C), .S00(N_185), .S01(N_187),
            .S1(N_140) );
csamuxb QL72 ( .A(N_200), .B(N_201), .Q(C15D), .S00(N_185), .S01(N_187),
            .S1(N_140) );
csamuxa QL73 ( .A(N_85), .Q(Q[18]), .S00(N_83), .S01(N_82), .S1(C15A) );
csamuxa QL74 ( .A(N_97), .Q(Q[20]), .S00(N_77), .S01(N_78), .S1(C15B) );
csamuxa QL75 ( .A(N_89), .Q(Q[24]), .S00(N_99), .S01(N_88), .S1(C15C) );
csamuxa QL76 ( .A(N_175), .Q(Q[10]), .S00(N_183), .S01(N_191), .S1(N_139) );
csamuxa QL77 ( .A(N_121), .Q(Q[6]), .S00(N_190), .S01(N_189), .S1(N_111) );
csamuxa QL78 ( .A(N_192), .Q(Q[12]), .S00(N_184), .S01(N_188), .S1(N_139) );
muxb2dx0 QL79 ( .A(N_74), .B(N_75), .C(N_74), .D(N_75), .Q(N_77), .R(N_2), .S(N_4),
             .T(N_83) );
muxb2dx0 QL80 ( .A(N_74), .B(N_75), .C(N_74), .D(N_75), .Q(N_78), .R(N_3), .S(N_76),
             .T(N_82) );
muxb2dx0 QL81 ( .A(N_15), .B(N_17), .C(N_18), .D(N_19), .Q(N_58), .R(N_59),
             .S(N_16), .T(N_57) );
muxb2dx0 QL82 ( .A(N_15), .B(N_17), .C(N_18), .D(N_19), .Q(N_62), .R(N_63),
             .S(N_20), .T(N_61) );
muxb2dx0 QL83 ( .A(N_176), .B(N_186), .C(N_176), .D(N_186), .Q(N_184), .R(N_185),
             .S(N_177), .T(N_183) );
muxb2dx0 QL84 ( .A(N_176), .B(N_186), .C(N_176), .D(N_186), .Q(N_188), .R(N_187),
             .S(N_178), .T(N_191) );
mux2x0 QL85 ( .A(N_54), .B(N_79), .Q(Q[17]), .S(C15A) );
mux2x0 QL86 ( .A(N_147), .B(N_148), .Q(Q[9]), .S(N_139) );
mux2dxx QL87 ( .A(N_92), .B(N_92), .C(N_90), .D(N_91), .Q(N_80), .R(N_81), .S(N_87) );
mux2dxx QL88 ( .A(N_48), .B(N_48), .C(N_50), .D(N_49), .Q(N_67), .R(N_68), .S(N_31) );
mux2dxx QL89 ( .A(N_48), .B(N_48), .C(N_50), .D(N_49), .Q(N_69), .R(N_70), .S(N_32) );
mux2dxx QL90 ( .A(N_64), .B(N_64), .C(N_65), .D(N_66), .Q(N_101), .R(N_102),
            .S(N_59) );
mux2dxx QL91 ( .A(N_64), .B(N_64), .C(N_65), .D(N_66), .Q(N_103), .R(N_104),
            .S(N_63) );
mux2dxx QL92 ( .A(N_92), .B(N_92), .C(N_90), .D(N_91), .Q(N_94), .R(N_93), .S(N_1) );
mux2dxx QL93 ( .A(N_199), .B(N_199), .C(N_160), .D(N_159), .Q(N_196), .R(N_182),
            .S(N_164) );
mux2dxx QL94 ( .A(N_199), .B(N_199), .C(N_160), .D(N_159), .Q(N_195), .R(N_197),
            .S(N_163) );
muxi2dx2 QL95 ( .A(N_5), .B(N_5), .C(N_7), .D(N_9), .Q(N_84), .R(N_75), .S(N_13) );
muxi2dx2 QL96 ( .A(N_6), .B(N_6), .C(N_8), .D(N_11), .Q(N_79), .R(N_76), .S(N_14) );
muxi2dx2 QL97 ( .A(N_21), .B(N_21), .C(N_23), .D(N_25), .Q(N_17), .R(N_19),
             .S(N_29) );
muxi2dx2 QL98 ( .A(N_22), .B(N_22), .C(N_24), .D(N_27), .Q(N_56), .R(N_20),
             .S(N_30) );
muxi2dx2 QL99 ( .A(N_33), .B(N_33), .C(N_34), .D(N_35), .Q(N_66), .R(N_32),
             .S(N_37) );
muxi2dx2 QL100 ( .A(N_38), .B(N_38), .C(N_40), .D(N_42), .Q(N_91), .R(N_98),
              .S(N_46) );
muxi2dx2 QL101 ( .A(N_39), .B(N_39), .C(N_41), .D(N_44), .Q(N_96), .R(N_87),
              .S(N_47) );
muxi2dx2 QL102 ( .A(N_145), .B(N_145), .C(N_144), .D(N_143), .Q(N_125), .R(N_122),
              .S(N_141) );
muxi2dx2 QL103 ( .A(N_149), .B(N_149), .C(N_151), .D(N_153), .Q(N_179), .R(N_186),
              .S(N_157) );
muxi2dx2 QL104 ( .A(N_150), .B(N_150), .C(N_152), .D(N_155), .Q(N_148), .R(N_178),
              .S(N_158) );
muxi2dx2 QL105 ( .A(N_165), .B(N_165), .C(N_167), .D(N_169), .Q(N_159), .R(N_161),
              .S(N_173) );
muxi2dx2 QL106 ( .A(N_166), .B(N_166), .C(N_168), .D(N_171), .Q(N_194), .R(N_164),
              .S(N_174) );
mux2dx2 QL107 ( .A(N_5), .B(N_5), .C(N_7), .D(N_9), .Q(N_86), .R(N_74), .S(N_10) );
mux2dx2 QL108 ( .A(N_6), .B(N_6), .C(N_8), .D(N_11), .Q(N_54), .R(N_4), .S(N_12) );
mux2dx2 QL109 ( .A(N_21), .B(N_21), .C(N_23), .D(N_25), .Q(N_15), .R(N_18),
             .S(N_26) );
mux2dx2 QL110 ( .A(N_22), .B(N_22), .C(N_24), .D(N_27), .Q(N_55), .R(N_16),
             .S(N_28) );
mux2dx2 QL111 ( .A(N_33), .B(N_33), .C(N_34), .D(N_35), .Q(N_65), .R(N_31),
             .S(N_36) );
mux2dx2 QL112 ( .A(N_38), .B(N_38), .C(N_40), .D(N_42), .Q(N_90), .R(N_100),
             .S(N_43) );
mux2dx2 QL113 ( .A(N_39), .B(N_39), .C(N_41), .D(N_44), .Q(N_95), .R(N_1), .S(N_45) );
mux2dx2 QL114 ( .A(N_57), .B(N_57), .C(N_61), .D(N_61), .Q(N_72), .R(N_71),
             .S(N_60) );
mux2dx2 QL115 ( .A(N_145), .B(N_145), .C(N_144), .D(N_143), .Q(N_126), .R(N_123),
             .S(N_142) );
mux2dx2 QL116 ( .A(N_149), .B(N_149), .C(N_151), .D(N_153), .Q(N_180), .R(N_176),
             .S(N_154) );
mux2dx2 QL117 ( .A(N_150), .B(N_150), .C(N_152), .D(N_155), .Q(N_147), .R(N_177),
             .S(N_156) );
mux2dx2 QL118 ( .A(N_165), .B(N_165), .C(N_167), .D(N_169), .Q(N_160), .R(N_162),
             .S(N_170) );
mux2dx2 QL119 ( .A(N_166), .B(N_166), .C(N_168), .D(N_171), .Q(N_193), .R(N_163),
             .S(N_172) );
mux2dx0 QL120 ( .A(N_67), .B(N_69), .C(N_68), .D(N_70), .Q(N_105), .R(N_106),
             .S(N_59) );
mux2dx0 QL121 ( .A(N_67), .B(N_69), .C(N_68), .D(N_70), .Q(N_107), .R(N_108),
             .S(N_63) );
mux2dx0 QL122 ( .A(N_162), .B(N_161), .C(N_162), .D(N_161), .Q(N_198), .R(N_200),
             .S(N_163) );
mux2dx0 QL123 ( .A(N_162), .B(N_161), .C(N_162), .D(N_161), .Q(N_181), .R(N_201),
             .S(N_164) );

endmodule // add32

`endif

`ifdef add16
`else
`define add16
module add16( A , B, Q );
 input [15:0] A;
 input [15:0] B;
 output [15:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;
wire N_15;
wire N_16;
wire N_17;
wire N_18;
wire N_19;
wire N_20;
wire N_21;
wire N_22;
wire N_23;
wire N_24;
wire N_25;
wire N_26;
wire N_27;
wire N_28;
wire N_29;
wire N_30;
wire N_31;
wire N_32;
wire N_33;
wire N_34;
wire N_35;
wire N_36;
wire N_37;
wire N_38;
wire N_39;
wire N_40;
wire N_41;
wire N_42;
wire N_43;
wire N_44;
wire N_45;
wire N_46;
wire N_47;
wire N_48;
wire N_49;
wire N_50;
wire N_51;
wire N_52;
wire N_53;
wire N_54;
wire N_55;
wire N_56;
wire N_57;
wire N_58;
wire N_59;
wire N_60;
wire N_61;
wire N_62;
wire N_63;
wire N_64;
wire N_65;
wire N_66;
wire N_67;
wire N_68;
wire N_69;
wire N_70;
wire N_71;
wire N_72;
wire N_73;
wire N_74;
wire N_75;
wire N_76;
wire N_77;
wire N_78;
wire N_79;
wire N_80;
wire N_81;
wire N_82;
wire N_83;

mux2dx2 QL1 ( .A(N_12), .B(N_12), .C(N_16), .D(N_23), .Q(N_61), .R(N_66), .S(N_24) );
mux2dx2 QL2 ( .A(N_11), .B(N_11), .C(N_15), .D(N_21), .Q(N_33), .R(N_4), .S(N_22) );
mux2dx2 QL3 ( .A(N_10), .B(N_10), .C(N_14), .D(N_19), .Q(N_3), .R(N_6), .S(N_20) );
mux2dx2 QL4 ( .A(N_9), .B(N_9), .C(N_13), .D(N_17), .Q(N_43), .R(N_2), .S(N_18) );
muxi2dx2 QL5 ( .A(N_12), .B(N_12), .C(N_16), .D(N_23), .Q(N_62), .R(N_67), .S(N_28) );
muxi2dx2 QL6 ( .A(N_11), .B(N_11), .C(N_15), .D(N_21), .Q(N_34), .R(N_8), .S(N_27) );
muxi2dx2 QL7 ( .A(N_10), .B(N_10), .C(N_14), .D(N_19), .Q(N_5), .R(N_7), .S(N_26) );
muxi2dx2 QL8 ( .A(N_9), .B(N_9), .C(N_13), .D(N_17), .Q(N_44), .R(N_29), .S(N_25) );
mux2dxx QL9 ( .A(N_1), .B(N_1), .C(N_80), .D(N_79), .Q(N_45), .R(N_46), .S(N_2) );
mux2dxx QL10 ( .A(N_1), .B(N_1), .C(N_80), .D(N_79), .Q(N_47), .R(N_48), .S(N_29) );
mux2x0 QL11 ( .A(N_33), .B(N_34), .Q(Q[9]), .S(N_31) );
mux2x0 QL12 ( .A(N_36), .B(N_40), .Q(Q[11]), .S(N_31) );
muxb2dx0 QL13 ( .A(N_3), .B(N_5), .C(N_6), .D(N_7), .Q(N_36), .R(N_37), .S(N_4),
             .T(N_35) );
muxb2dx0 QL14 ( .A(N_3), .B(N_5), .C(N_6), .D(N_7), .Q(N_40), .R(N_41), .S(N_8),
             .T(N_39) );
csamuxa QL15 ( .A(N_68), .Q(Q[6]), .S00(N_71), .S01(N_64), .S1(N_83) );
csamuxa QL16 ( .A(N_42), .Q(Q[12]), .S00(N_37), .S01(N_41), .S1(N_30) );
csamuxa QL17 ( .A(N_38), .Q(Q[10]), .S00(N_35), .S01(N_39), .S1(N_31) );
csamuxb QL18 ( .A(N_61), .B(N_62), .Q(Q[7]), .S00(N_71), .S01(N_64), .S1(N_83) );
csamuxb QL19 ( .A(N_43), .B(N_44), .Q(Q[13]), .S00(N_37), .S01(N_41), .S1(N_30) );
csamuxb QL20 ( .A(N_45), .B(N_47), .Q(Q[14]), .S00(N_37), .S01(N_41), .S1(N_30) );
csamuxb QL21 ( .A(N_46), .B(N_48), .Q(Q[15]), .S00(N_37), .S01(N_41), .S1(N_30) );
csamuxb QL22 ( .A(N_66), .B(N_67), .Q(N_31), .S00(N_63), .S01(N_65), .S1(N_69) );
csamuxb QL23 ( .A(N_66), .B(N_67), .Q(N_30), .S00(N_63), .S01(N_65), .S1(N_69) );
csamuxc QL24 ( .A(N_81), .B(N_82), .Q(N_69), .S00(N_50), .S01(N_51), .S1(N_53) );
csamuxd QL25 ( .A(N_49), .Q(Q[3]), .S00(N_50), .S01(N_51), .S1(N_74) );
csamuxd QL26 ( .A(N_60), .Q(Q[5]), .S00(N_70), .S01(N_72), .S1(N_83) );
mux4x6 QL27 ( .A(N_55), .B(N_55), .C(N_55), .D(N_55), .Q(Q[1]), .S0(N_52),
           .S1(B[1]) );
csalow QL28 ( .A0(A[0]), .A1(A[1]), .A1T(N_52), .B0(B[0]), .B1(B[1]), .C0(N_55),
           .C1(N_53) );
and2i2 QL29 ( .A(N_54), .B(N_55), .Q(Q[0]) );
nor2i0 QL30 ( .A(B[0]), .B(A[0]), .Q(N_54) );
muxb2dx2 QL31 ( .A(N_59), .B(N_58), .C(N_59), .D(N_58), .Q(N_71), .R(N_63),
             .S(N_56), .T(N_70) );
muxc2dx2 QL32 ( .A(N_59), .B(N_58), .C(N_59), .D(N_58), .Q(N_64), .R(N_65),
             .S(N_57), .T(N_72) );
buff QL33 ( .A(N_53), .Q(N_74) );
buff QL34 ( .A(N_69), .Q(N_83) );
csabita QL35 ( .A(A[4]), .B(B[4]), .C0(N_56), .C1(N_57), .S0(N_73) );
csabita QL36 ( .A(A[5]), .B(B[5]), .C0(N_59), .C1(N_58), .S0(N_60) );
csabita QL37 ( .A(A[6]), .B(B[6]), .C0(N_24), .C1(N_28), .S0(N_68) );
csabita QL38 ( .A(A[7]), .B(B[7]), .C0(N_16), .C1(N_23), .S0(N_12) );
csabita QL39 ( .A(A[8]), .B(B[8]), .C0(N_22), .C1(N_27), .S0(N_32) );
csabita QL40 ( .A(A[9]), .B(B[9]), .C0(N_15), .C1(N_21), .S0(N_11) );
csabita QL41 ( .A(A[10]), .B(B[10]), .C0(N_20), .C1(N_26), .S0(N_38) );
csabita QL42 ( .A(A[11]), .B(B[11]), .C0(N_14), .C1(N_19), .S0(N_10) );
csabita QL43 ( .A(A[12]), .B(B[12]), .C0(N_18), .C1(N_25), .S0(N_42) );
csabita QL44 ( .A(A[13]), .B(B[13]), .C0(N_13), .C1(N_17), .S0(N_9) );
csabita QL45 ( .A(A[14]), .B(B[14]), .C0(N_76), .C1(N_77), .S0(N_1) );
csabitb QL46 ( .A(A[2]), .B(B[2]), .C0(N_50), .C1(N_51), .S0(N_75) );
csabitb QL47 ( .A(A[3]), .B(B[3]), .C0(N_81), .C1(N_82), .S0(N_49) );
xor2p QL48 ( .A(N_74), .B(N_75), .Q(Q[2]) );
xor2p QL49 ( .A(N_83), .B(N_73), .Q(Q[4]) );
xor2p QL50 ( .A(N_31), .B(N_32), .Q(Q[8]) );
xor2p QL51 ( .A(A[15]), .B(B[15]), .Q(N_78) );
mux2dxy QL52 ( .A(N_76), .B(N_76), .C(N_77), .D(N_77), .Q(N_80), .R(N_79), .S(N_78) );

endmodule // add16

`endif

`ifdef accum8
`else
`define accum8
module accum8( A , CLK, CLR, Q );
 input [7:0] A;
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 output [7:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;
wire N_15;
wire N_16;
wire N_17;
wire N_18;
wire N_19;
wire N_20;
wire N_21;
wire N_22;
wire N_23;
wire N_24;
wire N_25;
wire N_26;
wire N_27;
wire N_28;
wire N_29;
wire N_30;
wire N_31;
wire N_32;
wire N_33;
wire N_34;
wire N_35;
wire N_36;
supply0 GND;

csamuxa QL1 ( .A(N_19), .Q(N_35), .S00(N_22), .S01(N_18), .S1(N_20) );
csamuxb QL2 ( .A(N_16), .B(N_17), .Q(N_36), .S00(N_22), .S01(N_18), .S1(N_20) );
csamuxc QL3 ( .A(N_27), .B(N_28), .Q(N_20), .S00(N_5), .S01(N_6), .S1(N_8) );
csamuxd QL4 ( .A(N_4), .Q(N_32), .S00(N_5), .S01(N_6), .S1(N_25) );
csamuxd QL5 ( .A(N_15), .Q(N_34), .S00(N_21), .S01(N_23), .S1(N_20) );
mux4x6 QL6 ( .A(N_10), .B(N_10), .C(N_10), .D(N_10), .Q(N_30), .S0(N_7), .S1(Q[1]) );
csalow QL7 ( .A0(A[0]), .A1(A[1]), .A1T(N_7), .B0(Q[0]), .B1(Q[1]), .C0(N_10),
          .C1(N_8) );
and2i2 QL8 ( .A(N_9), .B(N_10), .Q(N_29) );
nor2i0 QL9 ( .A(Q[0]), .B(A[0]), .Q(N_9) );
muxb2dx2 QL10 ( .A(N_14), .B(N_13), .C(GND), .D(GND), .Q(N_22), .S(N_11), .T(N_21) );
muxc2dx2 QL11 ( .A(N_14), .B(N_13), .C(GND), .D(GND), .Q(N_18), .S(N_12), .T(N_23) );
buff QL12 ( .A(N_8), .Q(N_25) );
csabita QL13 ( .A(A[4]), .B(Q[4]), .C0(N_11), .C1(N_12), .S0(N_24) );
csabita QL14 ( .A(A[5]), .B(Q[5]), .C0(N_14), .C1(N_13), .S0(N_15) );
csabita QL15 ( .A(A[6]), .B(Q[6]), .C0(N_2), .C1(N_3), .S0(N_19) );
csabita QL16 ( .A(A[7]), .B(Q[7]), .S0(N_1) );
csabitb QL17 ( .A(A[2]), .B(Q[2]), .C0(N_5), .C1(N_6), .S0(N_26) );
csabitb QL18 ( .A(A[3]), .B(Q[3]), .C0(N_27), .C1(N_28), .S0(N_4) );
xor2p QL19 ( .A(N_25), .B(N_26), .Q(N_31) );
xor2p QL20 ( .A(N_20), .B(N_24), .Q(N_33) );
dffc QL21 ( .CLK(CLK), .CLR(CLR), .D(N_29), .Q(Q[0]) );
dffc QL22 ( .CLK(CLK), .CLR(CLR), .D(N_30), .Q(Q[1]) );
dffc QL23 ( .CLK(CLK), .CLR(CLR), .D(N_31), .Q(Q[2]) );
dffc QL24 ( .CLK(CLK), .CLR(CLR), .D(N_32), .Q(Q[3]) );
dffc QL25 ( .CLK(CLK), .CLR(CLR), .D(N_33), .Q(Q[4]) );
dffc QL26 ( .CLK(CLK), .CLR(CLR), .D(N_34), .Q(Q[5]) );
dffc QL27 ( .CLK(CLK), .CLR(CLR), .D(N_35), .Q(Q[6]) );
dffc QL28 ( .CLK(CLK), .CLR(CLR), .D(N_36), .Q(Q[7]) );
mux2x2 QL29 ( .A(N_1), .B(N_1), .Q(N_16), .S(N_2) );
mux2x1 QL30 ( .A(N_1), .B(N_1), .Q(N_17), .S(N_3) );

endmodule // accum8

`endif

`ifdef accum4
`else
`define accum4
module accum4( A , CLK, CLR, Q );
 input [3:0] A;
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 output [3:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;

csamuxd QL1 ( .A(N_1), .Q(N_12), .S00(N_2), .S01(N_3), .S1(N_5) );
mux4x6 QL2 ( .A(N_7), .B(N_7), .C(N_7), .D(N_7), .Q(N_10), .S0(N_4), .S1(Q[1]) );
csalow QL3 ( .A0(A[0]), .A1(A[1]), .A1T(N_4), .B0(Q[0]), .B1(Q[1]), .C0(N_7),
          .C1(N_5) );
and2i2 QL4 ( .A(N_6), .B(N_7), .Q(N_9) );
nor2i0 QL5 ( .A(Q[0]), .B(A[0]), .Q(N_6) );
csabitb QL6 ( .A(A[2]), .B(Q[2]), .C0(N_2), .C1(N_3), .S0(N_8) );
csabitb QL7 ( .A(A[3]), .B(Q[3]), .S0(N_1) );
xor2p QL8 ( .A(N_5), .B(N_8), .Q(N_11) );
dffc QL9 ( .CLK(CLK), .CLR(CLR), .D(N_9), .Q(Q[0]) );
dffc QL10 ( .CLK(CLK), .CLR(CLR), .D(N_10), .Q(Q[1]) );
dffc QL11 ( .CLK(CLK), .CLR(CLR), .D(N_11), .Q(Q[2]) );
dffc QL12 ( .CLK(CLK), .CLR(CLR), .D(N_12), .Q(Q[3]) );

endmodule // accum4

`endif

`ifdef accum32
`else
`define accum32
module accum32( A , CLK, CLR, Q );
 input [31:0] A;
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 output [31:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;
wire N_15;
wire N_16;
wire N_17;
wire N_18;
wire N_19;
wire N_20;
wire N_21;
wire N_22;
wire N_23;
wire N_24;
wire N_25;
wire N_26;
wire N_27;
wire N_28;
wire N_29;
wire N_30;
wire N_31;
wire N_32;
wire N_33;
wire N_34;
wire N_35;
wire N_36;
wire N_37;
wire N_38;
wire N_39;
wire N_40;
wire N_41;
wire N_42;
wire N_43;
wire N_44;
wire N_45;
wire N_46;
wire N_47;
wire N_48;
wire N_49;
wire N_50;
wire N_51;
wire N_52;
wire N_53;
wire N_54;
wire N_55;
wire N_56;
wire N_57;
wire N_58;
wire N_59;
wire N_60;
wire N_61;
wire N_62;
wire N_63;
wire N_64;
wire N_65;
wire N_66;
wire N_67;
wire N_68;
wire N_69;
wire N_70;
wire N_71;
wire N_72;
wire N_73;
wire N_74;
wire N_75;
wire N_76;
wire N_77;
wire N_78;
wire N_79;
wire N_80;
wire N_81;
wire N_82;
wire N_83;
wire N_84;
wire N_85;
wire N_86;
wire N_87;
wire N_88;
wire N_89;
wire N_90;
wire N_91;
wire N_92;
wire N_93;
wire N_94;
wire N_95;
wire N_96;
wire N_97;
wire N_98;
wire N_99;
wire N_100;
wire N_101;
wire N_102;
wire N_103;
wire N_104;
wire N_105;
wire N_106;
wire N_107;
wire N_108;
wire N_109;
wire N_110;
wire N_111;
wire N_112;
wire N_113;
wire N_114;
wire N_115;
wire N_116;
wire N_117;
wire N_118;
wire N_119;
wire N_120;
wire N_121;
wire N_122;
wire N_123;
wire N_124;
wire N_125;
wire N_126;
wire N_127;
wire N_128;
wire N_129;
wire N_130;
wire N_131;
wire N_132;
wire N_133;
wire N_134;
wire N_135;
wire N_136;
wire N_137;
wire N_138;
wire N_139;
wire N_140;
wire N_141;
wire N_142;
wire N_143;
wire N_144;
wire N_145;
wire N_146;
wire N_147;
wire N_148;
wire N_149;
wire N_150;
wire N_151;
wire N_152;
wire N_153;
wire N_154;
wire N_155;
wire N_156;
wire N_157;
wire N_158;
wire N_159;
wire N_160;
wire N_161;
wire N_162;
wire N_163;
wire N_164;
wire N_165;
wire N_166;
wire N_167;
wire N_168;
wire N_169;
wire N_170;
wire N_171;
wire N_172;
wire N_173;
wire N_174;
wire N_175;
wire N_176;
wire N_177;
wire N_178;
wire N_179;
wire N_180;
wire N_181;
wire N_182;
wire N_183;
wire N_184;
wire N_185;
wire N_186;
wire N_187;
wire N_188;
wire N_189;
wire N_190;
wire N_191;
wire N_192;
wire N_193;
wire N_194;
wire N_195;
wire N_196;
wire N_197;
wire N_198;
wire N_199;
wire N_200;
wire N_201;
wire N_202;
wire N_203;
wire N_204;
wire N_205;
wire N_206;
wire N_207;
wire N_208;
wire N_209;
wire N_210;
wire N_211;
wire N_212;
wire N_213;
wire N_214;
wire N_215;
wire N_216;
wire N_217;
wire N_218;
wire N_219;
wire N_220;
wire N_221;
wire N_222;
wire C15A;
wire C15B;
wire N_223;
wire N_224;
wire N_225;
wire N_226;
wire N_227;
wire N_228;
wire N_229;
wire N_230;
wire C15C;
wire C15D;
wire N_231;
wire N_232;
wire N_233;

mux2dxy QL1 ( .A(N_52), .B(N_52), .C(N_53), .D(N_53), .Q(N_50), .R(N_49), .S(N_51) );
dffc QL2 ( .CLK(CLK), .CLR(CLR), .D(N_85), .Q(Q[17]) );
dffc QL3 ( .CLK(CLK), .CLR(CLR), .D(N_86), .Q(Q[16]) );
dffc QL4 ( .CLK(CLK), .CLR(CLR), .D(N_84), .Q(Q[18]) );
dffc QL5 ( .CLK(CLK), .CLR(CLR), .D(N_80), .Q(Q[23]) );
dffc QL6 ( .CLK(CLK), .CLR(CLR), .D(N_81), .Q(Q[22]) );
dffc QL7 ( .CLK(CLK), .CLR(CLR), .D(N_82), .Q(Q[21]) );
dffc QL8 ( .CLK(CLK), .CLR(CLR), .D(N_83), .Q(Q[20]) );
dffc QL9 ( .CLK(CLK), .CLR(CLR), .D(N_79), .Q(Q[25]) );
dffc QL10 ( .CLK(CLK), .CLR(CLR), .D(N_78), .Q(Q[26]) );
dffc QL11 ( .CLK(CLK), .CLR(CLR), .D(N_77), .Q(Q[27]) );
dffc QL12 ( .CLK(CLK), .CLR(CLR), .D(N_76), .Q(Q[28]) );
dffc QL13 ( .CLK(CLK), .CLR(CLR), .D(N_75), .Q(Q[29]) );
dffc QL14 ( .CLK(CLK), .CLR(CLR), .D(N_74), .Q(Q[30]) );
dffc QL15 ( .CLK(CLK), .CLR(CLR), .D(N_73), .Q(Q[31]) );
dffc QL16 ( .CLK(CLK), .CLR(CLR), .D(N_99), .Q(Q[19]) );
dffc QL17 ( .CLK(CLK), .CLR(CLR), .D(N_103), .Q(Q[24]) );
dffc QL18 ( .CLK(CLK), .CLR(CLR), .D(N_128), .Q(Q[7]) );
dffc QL19 ( .CLK(CLK), .CLR(CLR), .D(N_129), .Q(Q[6]) );
dffc QL20 ( .CLK(CLK), .CLR(CLR), .D(N_130), .Q(Q[5]) );
dffc QL21 ( .CLK(CLK), .CLR(CLR), .D(N_131), .Q(Q[4]) );
dffc QL22 ( .CLK(CLK), .CLR(CLR), .D(N_132), .Q(Q[3]) );
dffc QL23 ( .CLK(CLK), .CLR(CLR), .D(N_133), .Q(Q[2]) );
dffc QL24 ( .CLK(CLK), .CLR(CLR), .D(N_134), .Q(Q[1]) );
dffc QL25 ( .CLK(CLK), .CLR(CLR), .D(N_135), .Q(Q[0]) );
dffc QL26 ( .CLK(CLK), .CLR(CLR), .D(N_127), .Q(Q[10]) );
dffc QL27 ( .CLK(CLK), .CLR(CLR), .D(N_184), .Q(Q[9]) );
dffc QL28 ( .CLK(CLK), .CLR(CLR), .D(N_185), .Q(Q[8]) );
dffc QL29 ( .CLK(CLK), .CLR(CLR), .D(N_202), .Q(Q[15]) );
dffc QL30 ( .CLK(CLK), .CLR(CLR), .D(N_203), .Q(Q[14]) );
dffc QL31 ( .CLK(CLK), .CLR(CLR), .D(N_204), .Q(Q[13]) );
dffc QL32 ( .CLK(CLK), .CLR(CLR), .D(N_205), .Q(Q[12]) );
dffc QL33 ( .CLK(CLK), .CLR(CLR), .D(N_206), .Q(Q[11]) );
xor2p QL34 ( .A(A[31]), .B(Q[31]), .Q(N_51) );
xor2p QL35 ( .A(C15A), .B(N_87), .Q(N_86) );
xor2p QL36 ( .A(N_164), .B(N_171), .Q(N_185) );
xor2p QL37 ( .A(N_136), .B(N_141), .Q(N_131) );
xor2p QL38 ( .A(N_140), .B(N_139), .Q(N_133) );
csabitb QL39 ( .A(A[3]), .B(Q[3]), .C0(N_138), .C1(N_137), .S0(N_163) );
csabitb QL40 ( .A(A[2]), .B(Q[2]), .C0(N_162), .C1(N_161), .S0(N_139) );
csabita QL41 ( .A(A[18]), .B(Q[18]), .C0(N_10), .C1(N_13), .S0(N_100) );
csabita QL42 ( .A(A[19]), .B(Q[19]), .C0(N_7), .C1(N_9), .S0(N_5) );
csabita QL43 ( .A(A[20]), .B(Q[20]), .C0(N_45), .C1(N_47), .S0(N_113) );
csabita QL44 ( .A(A[21]), .B(Q[21]), .C0(N_41), .C1(N_44), .S0(N_39) );
csabita QL45 ( .A(A[22]), .B(Q[22]), .C0(N_43), .C1(N_46), .S0(N_108) );
csabita QL46 ( .A(A[23]), .B(Q[23]), .C0(N_40), .C1(N_42), .S0(N_38) );
csabita QL47 ( .A(A[24]), .B(Q[24]), .C0(N_28), .C1(N_30), .S0(N_105) );
csabita QL48 ( .A(A[25]), .B(Q[25]), .C0(N_24), .C1(N_27), .S0(N_22) );
csabita QL49 ( .A(A[26]), .B(Q[26]), .C0(N_26), .C1(N_29), .S0(N_60) );
csabita QL50 ( .A(A[27]), .B(Q[27]), .C0(N_23), .C1(N_25), .S0(N_21) );
csabita QL51 ( .A(A[28]), .B(Q[28]), .C0(N_36), .C1(N_37), .S0(N_64) );
csabita QL52 ( .A(A[29]), .B(Q[29]), .C0(N_34), .C1(N_35), .S0(N_33) );
csabita QL53 ( .A(A[30]), .B(Q[30]), .C0(N_52), .C1(N_53), .S0(N_48) );
csabita QL54 ( .A(A[17]), .B(Q[17]), .C0(N_8), .C1(N_11), .S0(N_6) );
csabita QL55 ( .A(A[16]), .B(Q[16]), .C0(N_12), .C1(N_14), .S0(N_87) );
csabita QL56 ( .A(A[14]), .B(Q[14]), .C0(N_197), .C1(N_200), .S0(N_231) );
csabita QL57 ( .A(A[13]), .B(Q[13]), .C0(N_195), .C1(N_198), .S0(N_193) );
csabita QL58 ( .A(A[12]), .B(Q[12]), .C0(N_199), .C1(N_201), .S0(N_224) );
csabita QL59 ( .A(A[11]), .B(Q[11]), .C0(N_176), .C1(N_178), .S0(N_174) );
csabita QL60 ( .A(A[10]), .B(Q[10]), .C0(N_179), .C1(N_182), .S0(N_207) );
csabita QL61 ( .A(A[9]), .B(Q[9]), .C0(N_177), .C1(N_180), .S0(N_175) );
csabita QL62 ( .A(A[8]), .B(Q[8]), .C0(N_181), .C1(N_183), .S0(N_171) );
csabita QL63 ( .A(A[7]), .B(Q[7]), .C0(N_169), .C1(N_168), .S0(N_170) );
csabita QL64 ( .A(A[6]), .B(Q[6]), .C0(N_167), .C1(N_166), .S0(N_146) );
csabita QL65 ( .A(A[5]), .B(Q[5]), .C0(N_153), .C1(N_154), .S0(N_152) );
csabita QL66 ( .A(A[4]), .B(Q[4]), .C0(N_156), .C1(N_155), .S0(N_141) );
csabita QL67 ( .A(A[15]), .B(Q[15]), .C0(N_194), .C1(N_196), .S0(N_192) );
buff QL68 ( .A(N_145), .Q(N_136) );
buff QL69 ( .A(N_159), .Q(N_140) );
muxc2dx2 QL70 ( .A(N_153), .B(N_154), .C(N_153), .D(N_154), .Q(N_221), .R(N_149),
             .S(N_155), .T(N_142) );
muxb2dx2 QL71 ( .A(N_153), .B(N_154), .C(N_153), .D(N_154), .Q(N_222), .R(N_143),
             .S(N_156), .T(N_144) );
nor2i0 QL72 ( .A(Q[0]), .B(A[0]), .Q(N_158) );
and2i2 QL73 ( .A(N_158), .B(N_157), .Q(N_135) );
csalow QL74 ( .A0(A[0]), .A1(A[1]), .A1T(N_160), .B0(Q[0]), .B1(Q[1]), .C0(N_157),
           .C1(N_159) );
mux4x6 QL75 ( .A(N_157), .B(N_157), .C(N_157), .D(N_157), .Q(N_134), .S0(N_160),
           .S1(Q[1]) );
csamuxd QL76 ( .A(N_152), .Q(N_130), .S00(N_144), .S01(N_142), .S1(N_136) );
csamuxd QL77 ( .A(N_163), .Q(N_132), .S00(N_162), .S01(N_161), .S1(N_140) );
csamuxc QL78 ( .A(N_138), .B(N_137), .Q(N_145), .S00(N_162), .S01(N_161),
            .S1(N_159) );
csamuxb QL79 ( .A(N_109), .B(N_95), .Q(N_80), .S00(N_91), .S01(N_92), .S1(C15B) );
csamuxb QL80 ( .A(N_110), .B(N_94), .Q(N_81), .S00(N_91), .S01(N_92), .S1(C15B) );
csamuxb QL81 ( .A(N_111), .B(N_112), .Q(N_82), .S00(N_91), .S01(N_92), .S1(C15B) );
csamuxb QL82 ( .A(N_55), .B(N_56), .Q(N_79), .S00(N_115), .S01(N_104), .S1(C15C) );
csamuxb QL83 ( .A(N_72), .B(N_71), .Q(N_78), .S00(N_115), .S01(N_104), .S1(C15C) );
csamuxb QL84 ( .A(N_58), .B(N_62), .Q(N_77), .S00(N_115), .S01(N_104), .S1(C15C) );
csamuxb QL85 ( .A(N_117), .B(N_119), .Q(N_76), .S00(N_126), .S01(N_125), .S1(C15D) );
csamuxb QL86 ( .A(N_118), .B(N_120), .Q(N_75), .S00(N_126), .S01(N_125), .S1(C15D) );
csamuxb QL87 ( .A(N_121), .B(N_123), .Q(N_74), .S00(N_126), .S01(N_125), .S1(C15D) );
csamuxb QL88 ( .A(N_122), .B(N_124), .Q(N_73), .S00(N_126), .S01(N_125), .S1(C15D) );
csamuxb QL89 ( .A(N_101), .B(N_98), .Q(N_99), .S00(N_97), .S01(N_96), .S1(C15A) );
csamuxb QL90 ( .A(N_116), .B(N_114), .Q(N_104), .S00(N_1), .S01(N_102), .S1(N_3) );
csamuxb QL91 ( .A(N_116), .B(N_114), .Q(N_115), .S00(N_1), .S01(N_102), .S1(N_2) );
csamuxb QL92 ( .A(N_116), .B(N_114), .Q(N_126), .S00(N_1), .S01(N_102), .S1(N_2) );
csamuxb QL93 ( .A(N_116), .B(N_114), .Q(N_125), .S00(N_1), .S01(N_102), .S1(N_3) );
csamuxb QL94 ( .A(N_148), .B(N_147), .Q(N_165), .S00(N_143), .S01(N_149),
            .S1(N_145) );
csamuxb QL95 ( .A(N_148), .B(N_147), .Q(N_164), .S00(N_222), .S01(N_221),
            .S1(N_145) );
csamuxb QL96 ( .A(N_225), .B(N_226), .Q(N_204), .S00(N_216), .S01(N_220),
            .S1(N_164) );
csamuxb QL97 ( .A(N_151), .B(N_150), .Q(N_128), .S00(N_222), .S01(N_221),
            .S1(N_136) );
csamuxb QL98 ( .A(N_230), .B(N_213), .Q(C15A), .S00(N_217), .S01(N_219),
            .S1(N_165) );
csamuxb QL99 ( .A(N_229), .B(N_214), .Q(N_202), .S00(N_216), .S01(N_220),
            .S1(N_164) );
csamuxb QL100 ( .A(N_227), .B(N_228), .Q(N_203), .S00(N_216), .S01(N_220),
             .S1(N_164) );
csamuxb QL101 ( .A(N_212), .B(N_211), .Q(N_206), .S00(N_215), .S01(N_223),
             .S1(N_164) );
csamuxb QL102 ( .A(N_230), .B(N_213), .Q(C15B), .S00(N_217), .S01(N_219),
             .S1(N_165) );
csamuxb QL103 ( .A(N_232), .B(N_233), .Q(C15C), .S00(N_217), .S01(N_219),
             .S1(N_165) );
csamuxb QL104 ( .A(N_232), .B(N_233), .Q(C15D), .S00(N_217), .S01(N_219),
             .S1(N_165) );
csamuxa QL105 ( .A(N_100), .Q(N_84), .S00(N_97), .S01(N_96), .S1(C15A) );
csamuxa QL106 ( .A(N_113), .Q(N_83), .S00(N_91), .S01(N_92), .S1(C15B) );
csamuxa QL107 ( .A(N_105), .Q(N_103), .S00(N_115), .S01(N_104), .S1(C15C) );
csamuxa QL108 ( .A(N_207), .Q(N_127), .S00(N_215), .S01(N_223), .S1(N_164) );
csamuxa QL109 ( .A(N_146), .Q(N_129), .S00(N_222), .S01(N_221), .S1(N_136) );
csamuxa QL110 ( .A(N_224), .Q(N_205), .S00(N_216), .S01(N_220), .S1(N_164) );
muxb2dx0 QL111 ( .A(N_88), .B(N_89), .C(N_88), .D(N_89), .Q(N_91), .R(N_2), .S(N_4),
              .T(N_97) );
muxb2dx0 QL112 ( .A(N_88), .B(N_89), .C(N_88), .D(N_89), .Q(N_92), .R(N_3),
              .S(N_90), .T(N_96) );
muxb2dx0 QL113 ( .A(N_15), .B(N_17), .C(N_18), .D(N_19), .Q(N_58), .R(N_59),
              .S(N_16), .T(N_57) );
muxb2dx0 QL114 ( .A(N_15), .B(N_17), .C(N_18), .D(N_19), .Q(N_62), .R(N_63),
              .S(N_20), .T(N_61) );
muxb2dx0 QL115 ( .A(N_208), .B(N_218), .C(N_208), .D(N_218), .Q(N_216), .R(N_217),
              .S(N_209), .T(N_215) );
muxb2dx0 QL116 ( .A(N_208), .B(N_218), .C(N_208), .D(N_218), .Q(N_220), .R(N_219),
              .S(N_210), .T(N_223) );
mux2x0 QL117 ( .A(N_54), .B(N_93), .Q(N_85), .S(C15A) );
mux2x0 QL118 ( .A(N_172), .B(N_173), .Q(N_184), .S(N_164) );
mux2dxx QL119 ( .A(N_108), .B(N_108), .C(N_106), .D(N_107), .Q(N_94), .R(N_95),
             .S(N_102) );
mux2dxx QL120 ( .A(N_48), .B(N_48), .C(N_50), .D(N_49), .Q(N_67), .R(N_68),
             .S(N_31) );
mux2dxx QL121 ( .A(N_48), .B(N_48), .C(N_50), .D(N_49), .Q(N_69), .R(N_70),
             .S(N_32) );
mux2dxx QL122 ( .A(N_64), .B(N_64), .C(N_65), .D(N_66), .Q(N_117), .R(N_118),
             .S(N_59) );
mux2dxx QL123 ( .A(N_64), .B(N_64), .C(N_65), .D(N_66), .Q(N_119), .R(N_120),
             .S(N_63) );
mux2dxx QL124 ( .A(N_108), .B(N_108), .C(N_106), .D(N_107), .Q(N_110), .R(N_109),
             .S(N_1) );
mux2dxx QL125 ( .A(N_231), .B(N_231), .C(N_187), .D(N_186), .Q(N_228), .R(N_214),
             .S(N_191) );
mux2dxx QL126 ( .A(N_231), .B(N_231), .C(N_187), .D(N_186), .Q(N_227), .R(N_229),
             .S(N_190) );
muxi2dx2 QL127 ( .A(N_5), .B(N_5), .C(N_7), .D(N_9), .Q(N_98), .R(N_89), .S(N_13) );
muxi2dx2 QL128 ( .A(N_6), .B(N_6), .C(N_8), .D(N_11), .Q(N_93), .R(N_90), .S(N_14) );
muxi2dx2 QL129 ( .A(N_21), .B(N_21), .C(N_23), .D(N_25), .Q(N_17), .R(N_19),
              .S(N_29) );
muxi2dx2 QL130 ( .A(N_22), .B(N_22), .C(N_24), .D(N_27), .Q(N_56), .R(N_20),
              .S(N_30) );
muxi2dx2 QL131 ( .A(N_33), .B(N_33), .C(N_34), .D(N_35), .Q(N_66), .R(N_32),
              .S(N_37) );
muxi2dx2 QL132 ( .A(N_38), .B(N_38), .C(N_40), .D(N_42), .Q(N_107), .R(N_114),
              .S(N_46) );
muxi2dx2 QL133 ( .A(N_39), .B(N_39), .C(N_41), .D(N_44), .Q(N_112), .R(N_102),
              .S(N_47) );
muxi2dx2 QL134 ( .A(N_170), .B(N_170), .C(N_169), .D(N_168), .Q(N_150), .R(N_147),
              .S(N_166) );
muxi2dx2 QL135 ( .A(N_174), .B(N_174), .C(N_176), .D(N_178), .Q(N_211), .R(N_218),
              .S(N_182) );
muxi2dx2 QL136 ( .A(N_175), .B(N_175), .C(N_177), .D(N_180), .Q(N_173), .R(N_210),
              .S(N_183) );
muxi2dx2 QL137 ( .A(N_192), .B(N_192), .C(N_194), .D(N_196), .Q(N_186), .R(N_188),
              .S(N_200) );
muxi2dx2 QL138 ( .A(N_193), .B(N_193), .C(N_195), .D(N_198), .Q(N_226), .R(N_191),
              .S(N_201) );
mux2dx2 QL139 ( .A(N_5), .B(N_5), .C(N_7), .D(N_9), .Q(N_101), .R(N_88), .S(N_10) );
mux2dx2 QL140 ( .A(N_6), .B(N_6), .C(N_8), .D(N_11), .Q(N_54), .R(N_4), .S(N_12) );
mux2dx2 QL141 ( .A(N_21), .B(N_21), .C(N_23), .D(N_25), .Q(N_15), .R(N_18),
             .S(N_26) );
mux2dx2 QL142 ( .A(N_22), .B(N_22), .C(N_24), .D(N_27), .Q(N_55), .R(N_16),
             .S(N_28) );
mux2dx2 QL143 ( .A(N_33), .B(N_33), .C(N_34), .D(N_35), .Q(N_65), .R(N_31),
             .S(N_36) );
mux2dx2 QL144 ( .A(N_38), .B(N_38), .C(N_40), .D(N_42), .Q(N_106), .R(N_116),
             .S(N_43) );
mux2dx2 QL145 ( .A(N_39), .B(N_39), .C(N_41), .D(N_44), .Q(N_111), .R(N_1),
             .S(N_45) );
mux2dx2 QL146 ( .A(N_57), .B(N_57), .C(N_61), .D(N_61), .Q(N_72), .R(N_71),
             .S(N_60) );
mux2dx2 QL147 ( .A(N_170), .B(N_170), .C(N_169), .D(N_168), .Q(N_151), .R(N_148),
             .S(N_167) );
mux2dx2 QL148 ( .A(N_174), .B(N_174), .C(N_176), .D(N_178), .Q(N_212), .R(N_208),
             .S(N_179) );
mux2dx2 QL149 ( .A(N_175), .B(N_175), .C(N_177), .D(N_180), .Q(N_172), .R(N_209),
             .S(N_181) );
mux2dx2 QL150 ( .A(N_192), .B(N_192), .C(N_194), .D(N_196), .Q(N_187), .R(N_189),
             .S(N_197) );
mux2dx2 QL151 ( .A(N_193), .B(N_193), .C(N_195), .D(N_198), .Q(N_225), .R(N_190),
             .S(N_199) );
mux2dx0 QL152 ( .A(N_67), .B(N_69), .C(N_68), .D(N_70), .Q(N_121), .R(N_122),
             .S(N_59) );
mux2dx0 QL153 ( .A(N_67), .B(N_69), .C(N_68), .D(N_70), .Q(N_123), .R(N_124),
             .S(N_63) );
mux2dx0 QL154 ( .A(N_189), .B(N_188), .C(N_189), .D(N_188), .Q(N_230), .R(N_232),
             .S(N_190) );
mux2dx0 QL155 ( .A(N_189), .B(N_188), .C(N_189), .D(N_188), .Q(N_213), .R(N_233),
             .S(N_191) );

endmodule // accum32

`endif

`ifdef accum16
`else
`define accum16
module accum16( A , CLK, CLR, Q );
 input [15:0] A;
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 output [15:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;
wire N_12;
wire N_13;
wire N_14;
wire N_15;
wire N_16;
wire N_17;
wire N_18;
wire N_19;
wire N_20;
wire N_21;
wire N_22;
wire N_23;
wire N_24;
wire N_25;
wire N_26;
wire N_27;
wire N_28;
wire N_29;
wire N_30;
wire N_31;
wire N_32;
wire N_33;
wire N_34;
wire N_35;
wire N_36;
wire N_37;
wire N_38;
wire N_39;
wire N_40;
wire N_41;
wire N_42;
wire N_43;
wire N_44;
wire N_45;
wire N_46;
wire N_47;
wire N_48;
wire N_49;
wire N_50;
wire N_51;
wire N_52;
wire N_53;
wire N_54;
wire N_55;
wire N_56;
wire N_57;
wire N_58;
wire N_59;
wire N_60;
wire N_61;
wire N_62;
wire N_63;
wire N_64;
wire N_65;
wire N_66;
wire N_67;
wire N_68;
wire N_69;
wire N_70;
wire N_71;
wire N_72;
wire N_73;
wire N_74;
wire N_75;
wire N_76;
wire N_77;
wire N_78;
wire N_79;
wire N_80;
wire N_81;
wire N_82;
wire N_83;
wire N_84;
wire N_85;
wire N_86;
wire N_87;
wire N_88;
wire N_89;
wire N_90;
wire N_91;
wire N_92;
wire N_93;
wire N_94;
wire N_95;
wire N_96;
wire N_97;
wire N_98;
wire N_99;

mux2dx2 QL1 ( .A(N_12), .B(N_12), .C(N_16), .D(N_23), .Q(N_61), .R(N_66), .S(N_24) );
mux2dx2 QL2 ( .A(N_11), .B(N_11), .C(N_15), .D(N_21), .Q(N_33), .R(N_4), .S(N_22) );
mux2dx2 QL3 ( .A(N_10), .B(N_10), .C(N_14), .D(N_19), .Q(N_3), .R(N_6), .S(N_20) );
mux2dx2 QL4 ( .A(N_9), .B(N_9), .C(N_13), .D(N_17), .Q(N_43), .R(N_2), .S(N_18) );
muxi2dx2 QL5 ( .A(N_12), .B(N_12), .C(N_16), .D(N_23), .Q(N_62), .R(N_67), .S(N_28) );
muxi2dx2 QL6 ( .A(N_11), .B(N_11), .C(N_15), .D(N_21), .Q(N_34), .R(N_8), .S(N_27) );
muxi2dx2 QL7 ( .A(N_10), .B(N_10), .C(N_14), .D(N_19), .Q(N_5), .R(N_7), .S(N_26) );
muxi2dx2 QL8 ( .A(N_9), .B(N_9), .C(N_13), .D(N_17), .Q(N_44), .R(N_29), .S(N_25) );
mux2dxx QL9 ( .A(N_1), .B(N_1), .C(N_80), .D(N_79), .Q(N_45), .R(N_46), .S(N_2) );
mux2dxx QL10 ( .A(N_1), .B(N_1), .C(N_80), .D(N_79), .Q(N_47), .R(N_48), .S(N_29) );
mux2x0 QL11 ( .A(N_33), .B(N_34), .Q(N_93), .S(N_31) );
mux2x0 QL12 ( .A(N_36), .B(N_40), .Q(N_94), .S(N_31) );
muxb2dx0 QL13 ( .A(N_3), .B(N_5), .C(N_6), .D(N_7), .Q(N_36), .R(N_37), .S(N_4),
             .T(N_35) );
muxb2dx0 QL14 ( .A(N_3), .B(N_5), .C(N_6), .D(N_7), .Q(N_40), .R(N_41), .S(N_8),
             .T(N_39) );
csamuxa QL15 ( .A(N_68), .Q(N_90), .S00(N_71), .S01(N_64), .S1(N_83) );
csamuxa QL16 ( .A(N_42), .Q(N_95), .S00(N_37), .S01(N_41), .S1(N_30) );
csamuxa QL17 ( .A(N_38), .Q(N_99), .S00(N_35), .S01(N_39), .S1(N_31) );
csamuxb QL18 ( .A(N_61), .B(N_62), .Q(N_91), .S00(N_71), .S01(N_64), .S1(N_83) );
csamuxb QL19 ( .A(N_43), .B(N_44), .Q(N_96), .S00(N_37), .S01(N_41), .S1(N_30) );
csamuxb QL20 ( .A(N_45), .B(N_47), .Q(N_97), .S00(N_37), .S01(N_41), .S1(N_30) );
csamuxb QL21 ( .A(N_46), .B(N_48), .Q(N_98), .S00(N_37), .S01(N_41), .S1(N_30) );
csamuxb QL22 ( .A(N_66), .B(N_67), .Q(N_31), .S00(N_63), .S01(N_65), .S1(N_69) );
csamuxb QL23 ( .A(N_66), .B(N_67), .Q(N_30), .S00(N_63), .S01(N_65), .S1(N_69) );
csamuxc QL24 ( .A(N_81), .B(N_82), .Q(N_69), .S00(N_50), .S01(N_51), .S1(N_53) );
csamuxd QL25 ( .A(N_49), .Q(N_87), .S00(N_50), .S01(N_51), .S1(N_74) );
csamuxd QL26 ( .A(N_60), .Q(N_89), .S00(N_70), .S01(N_72), .S1(N_83) );
mux4x6 QL27 ( .A(N_55), .B(N_55), .C(N_55), .D(N_55), .Q(N_85), .S0(N_52),
           .S1(Q[1]) );
csalow QL28 ( .A0(A[0]), .A1(A[1]), .A1T(N_52), .B0(Q[0]), .B1(Q[1]), .C0(N_55),
           .C1(N_53) );
and2i2 QL29 ( .A(N_54), .B(N_55), .Q(N_84) );
nor2i0 QL30 ( .A(Q[0]), .B(A[0]), .Q(N_54) );
muxb2dx2 QL31 ( .A(N_59), .B(N_58), .C(N_59), .D(N_58), .Q(N_71), .R(N_63),
             .S(N_56), .T(N_70) );
muxc2dx2 QL32 ( .A(N_59), .B(N_58), .C(N_59), .D(N_58), .Q(N_64), .R(N_65),
             .S(N_57), .T(N_72) );
buff QL33 ( .A(N_53), .Q(N_74) );
buff QL34 ( .A(N_69), .Q(N_83) );
csabita QL35 ( .A(A[4]), .B(Q[4]), .C0(N_56), .C1(N_57), .S0(N_73) );
csabita QL36 ( .A(A[5]), .B(Q[5]), .C0(N_59), .C1(N_58), .S0(N_60) );
csabita QL37 ( .A(A[6]), .B(Q[6]), .C0(N_24), .C1(N_28), .S0(N_68) );
csabita QL38 ( .A(A[7]), .B(Q[7]), .C0(N_16), .C1(N_23), .S0(N_12) );
csabita QL39 ( .A(A[8]), .B(Q[8]), .C0(N_22), .C1(N_27), .S0(N_32) );
csabita QL40 ( .A(A[9]), .B(Q[9]), .C0(N_15), .C1(N_21), .S0(N_11) );
csabita QL41 ( .A(A[10]), .B(Q[10]), .C0(N_20), .C1(N_26), .S0(N_38) );
csabita QL42 ( .A(A[11]), .B(Q[11]), .C0(N_14), .C1(N_19), .S0(N_10) );
csabita QL43 ( .A(A[12]), .B(Q[12]), .C0(N_18), .C1(N_25), .S0(N_42) );
csabita QL44 ( .A(A[13]), .B(Q[13]), .C0(N_13), .C1(N_17), .S0(N_9) );
csabita QL45 ( .A(A[14]), .B(Q[14]), .C0(N_76), .C1(N_77), .S0(N_1) );
csabitb QL46 ( .A(A[2]), .B(Q[2]), .C0(N_50), .C1(N_51), .S0(N_75) );
csabitb QL47 ( .A(A[3]), .B(Q[3]), .C0(N_81), .C1(N_82), .S0(N_49) );
xor2p QL48 ( .A(N_74), .B(N_75), .Q(N_86) );
xor2p QL49 ( .A(N_83), .B(N_73), .Q(N_88) );
xor2p QL50 ( .A(N_31), .B(N_32), .Q(N_92) );
xor2p QL51 ( .A(A[15]), .B(Q[15]), .Q(N_78) );
dffc QL52 ( .CLK(CLK), .CLR(CLR), .D(N_84), .Q(Q[0]) );
dffc QL53 ( .CLK(CLK), .CLR(CLR), .D(N_85), .Q(Q[1]) );
dffc QL54 ( .CLK(CLK), .CLR(CLR), .D(N_86), .Q(Q[2]) );
dffc QL55 ( .CLK(CLK), .CLR(CLR), .D(N_87), .Q(Q[3]) );
dffc QL56 ( .CLK(CLK), .CLR(CLR), .D(N_88), .Q(Q[4]) );
dffc QL57 ( .CLK(CLK), .CLR(CLR), .D(N_89), .Q(Q[5]) );
dffc QL58 ( .CLK(CLK), .CLR(CLR), .D(N_90), .Q(Q[6]) );
dffc QL59 ( .CLK(CLK), .CLR(CLR), .D(N_91), .Q(Q[7]) );
dffc QL60 ( .CLK(CLK), .CLR(CLR), .D(N_92), .Q(Q[8]) );
dffc QL61 ( .CLK(CLK), .CLR(CLR), .D(N_93), .Q(Q[9]) );
dffc QL62 ( .CLK(CLK), .CLR(CLR), .D(N_99), .Q(Q[10]) );
dffc QL63 ( .CLK(CLK), .CLR(CLR), .D(N_94), .Q(Q[11]) );
dffc QL64 ( .CLK(CLK), .CLR(CLR), .D(N_95), .Q(Q[12]) );
dffc QL65 ( .CLK(CLK), .CLR(CLR), .D(N_96), .Q(Q[13]) );
dffc QL66 ( .CLK(CLK), .CLR(CLR), .D(N_97), .Q(Q[14]) );
dffc QL67 ( .CLK(CLK), .CLR(CLR), .D(N_98), .Q(Q[15]) );
mux2dxy QL68 ( .A(N_76), .B(N_76), .C(N_77), .D(N_77), .Q(N_80), .R(N_79), .S(N_78) );

endmodule // accum16

`endif

`ifdef and14i7
`else
`define and14i7
module and14i7( A , B, C, D, E, F, G, H, I, J, K, L, M, N, Q );
input A, B, C, D, E, F, G, H, I, J, K, L, M, N;
output Q;
parameter syn_macro = 1, ql_pack = 1;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(A), .A2(H), .A3(B), .A4(I), .A5(C), .A6(J), .AZ(N_2) );
frag_f I_1 ( .F1(E), .F2(L), .F3(F), .F4(M), .F5(G), .F6(N), .FZ(N_1) );
frag_m QL3 ( .B1(GND), .B2(VCC), .C1(GND), .C2(VCC), .D1(GND), .D2(VCC), .E1(D),
          .E2(K), .NS(N_1), .OS(N_2), .OZ(Q) );

endmodule // and14i7

`endif

`ifdef upflct4a
`else
`define upflct4a
module upflct4a( CLK , CLR, D, LOAD, Q, RCO );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:3] D;
input LOAD;
 output [0:3] Q;
output RCO;
supply0 GND;
supply1 VCC;

upflbit QL5 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(Q[0]), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
upflbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(Q[1]), .Q0(Q[0]), .Q1(VCC), .Q2(VCC) );
upflbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(VCC) );
upflbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
nand2i0 QL1 ( .A(Q[2]), .B(Q[3]), .Q(RCO) );

endmodule // upflct4a

`endif

`ifdef upflct4b
`else
`define upflct4b
module upflct4b( CLK , CLR, D, ENP, ENT, LOAD, Q, RCO );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:3] D;
input ENP, ENT, LOAD;
 output [0:3] Q;
output RCO;
supply1 VCC;

upflbit QL5 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[0]), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
upflbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[1]), .Q0(Q[0]), .Q1(VCC), .Q2(VCC) );
upflbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(VCC) );
upflbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
nand5i1 QL1 ( .A(Q[0]), .B(Q[1]), .C(Q[2]), .D(Q[3]), .E(ENT), .Q(RCO) );

endmodule // upflct4b

`endif

`ifdef upflct4c
`else
`define upflct4c
module upflct4c( CLK , CLR, D, ENP, ENT, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:3] D;
input ENP, ENT, LOAD;
 output [0:3] Q;
supply1 VCC;

upflbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[0]), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
upflbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[1]), .Q0(Q[0]), .Q1(VCC), .Q2(VCC) );
upflbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(VCC) );
upflbit QL1 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );

endmodule // upflct4c

`endif

`ifdef upflcar2
`else
`define upflcar2
module upflcar2( CLK , CLR, D, LOAD, ACO1, ACO2 );
output ACO1, ACO2;
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:1] D;
input LOAD;
supply0 GND;
supply1 VCC;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;

and3i1 QL10 ( .A(D[0]), .B(D[1]), .C(LOAD), .Q(N_7) );
and3i1 QL9 ( .A(LOAD), .B(N_4), .C(N_3), .Q(N_5) );
and3i1 QL8 ( .A(D[0]), .B(D[1]), .C(LOAD), .Q(N_8) );
and3i1 QL7 ( .A(LOAD), .B(N_4), .C(N_3), .Q(N_6) );
mux4x0 QL6 ( .A(VCC), .B(GND), .C(GND), .D(VCC), .Q(N_1), .S0(N_5), .S1(N_7) );
mux4x0 QL5 ( .A(VCC), .B(GND), .C(GND), .D(VCC), .Q(N_2), .S0(N_6), .S1(N_8) );
upflbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(N_4), .Q0(N_3), .Q1(VCC), .Q2(VCC) );
upflbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(N_3), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
dffp QL2 ( .CLK(CLK), .D(N_2), .PRE(CLR), .Q(ACO2) );
dffp QL1 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO1) );

endmodule // upflcar2

`endif

`ifdef upflcar3
`else
`define upflcar3
module upflcar3( CLK , CLR, D, LOAD, ACO1, ACO2, ACO3 );
output ACO1, ACO2, ACO3;
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:1] D;
input LOAD;
supply1 VCC;
supply0 GND;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;

and3i1 QL14 ( .A(D[0]), .B(D[1]), .C(LOAD), .Q(N_9) );
and3i1 QL13 ( .A(LOAD), .B(N_5), .C(N_4), .Q(N_6) );
and3i1 QL12 ( .A(D[0]), .B(D[1]), .C(LOAD), .Q(N_10) );
and3i1 QL11 ( .A(LOAD), .B(N_5), .C(N_4), .Q(N_7) );
and3i1 QL10 ( .A(LOAD), .B(N_5), .C(N_4), .Q(N_8) );
and3i1 QL9 ( .A(D[0]), .B(D[1]), .C(LOAD), .Q(N_11) );
mux4x0 QL8 ( .A(VCC), .B(GND), .C(GND), .D(VCC), .Q(N_1), .S0(N_6), .S1(N_9) );
mux4x0 QL7 ( .A(VCC), .B(GND), .C(GND), .D(VCC), .Q(N_2), .S0(N_7), .S1(N_10) );
mux4x0 QL6 ( .A(VCC), .B(GND), .C(GND), .D(VCC), .Q(N_3), .S0(N_8), .S1(N_11) );
upflbit QL5 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(N_5), .Q0(N_4), .Q1(VCC), .Q2(VCC) );
upflbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(N_4), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
dffp QL3 ( .CLK(CLK), .D(N_3), .PRE(CLR), .Q(ACO3) );
dffp QL2 ( .CLK(CLK), .D(N_2), .PRE(CLR), .Q(ACO2) );
dffp QL1 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO1) );

endmodule // upflcar3

`endif

`ifdef upfxcar1
`else
`define upfxcar1
module upfxcar1( CLK , CLR, D, ENG, LOAD, Q, ACO1 );
output ACO1;
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:1] D;
input ENG, LOAD;
 input [0:1] Q;
wire N_1;
wire N_2;
wire N_3;

mux4x7 QL4 ( .A(N_2), .B(N_2), .C(N_3), .D(ACO1), .Q(N_1), .S0(ENG), .S1(LOAD) );
and2i1 QL3 ( .A(Q[1]), .B(Q[0]), .Q(N_3) );
and2i0 QL2 ( .A(D[0]), .B(D[1]), .Q(N_2) );
dffp QL1 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO1) );

endmodule // upfxcar1

`endif

`ifdef upfxct4c
`else
`define upfxct4c
module upfxct4c( CLK , CLR, D, ENG, ENP, ENT, LOAD, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:3] D;
input ENG, ENP, ENT, LOAD;
 output [0:3] Q;
supply1 VCC;

upfxbit QL1 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
upfxbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(VCC) );
upfxbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[1]), .Q0(Q[0]), .Q1(VCC), .Q2(VCC) );
upfxbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[0]), .Q0(VCC), .Q1(VCC), .Q2(VCC) );

endmodule // upfxct4c

`endif

`ifdef upfxct4a
`else
`define upfxct4a
module upfxct4a( CLK , CLR, D, ENG, LOAD, Q, RCO );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:3] D;
input ENG, LOAD;
 output [0:3] Q;
output RCO;
supply0 GND;
supply1 VCC;

nand2i0 QL1 ( .A(Q[2]), .B(Q[3]), .Q(RCO) );
upfxbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENG(ENG), .ENP(GND), .ENT(GND),
           .LOAD(LOAD), .Q(Q[0]), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
upfxbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENG(ENG), .ENP(GND), .ENT(GND),
           .LOAD(LOAD), .Q(Q[1]), .Q0(Q[0]), .Q1(VCC), .Q2(VCC) );
upfxbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENG(ENG), .ENP(GND), .ENT(GND),
           .LOAD(LOAD), .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(VCC) );
upfxbit QL5 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENG(ENG), .ENP(GND), .ENT(GND),
           .LOAD(LOAD), .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );

endmodule // upfxct4a

`endif

`ifdef upfxcar3
`else
`define upfxcar3
module upfxcar3( CLK , CLR, D, ENG, LOAD, Q, ACO1, ACO2, ACO3 );
output ACO1, ACO2, ACO3;
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:1] D;
input ENG, LOAD;
 input [0:1] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;

mux4x7 QL8 ( .A(N_4), .B(N_4), .C(N_5), .D(ACO3), .Q(N_1), .S0(ENG), .S1(LOAD) );
mux4x7 QL7 ( .A(N_4), .B(N_4), .C(N_5), .D(ACO2), .Q(N_2), .S0(ENG), .S1(LOAD) );
mux4x7 QL6 ( .A(N_4), .B(N_4), .C(N_5), .D(ACO1), .Q(N_3), .S0(ENG), .S1(LOAD) );
and2i1 QL5 ( .A(Q[1]), .B(Q[0]), .Q(N_5) );
and2i0 QL4 ( .A(D[0]), .B(D[1]), .Q(N_4) );
dffp QL3 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO3) );
dffp QL2 ( .CLK(CLK), .D(N_2), .PRE(CLR), .Q(ACO2) );
dffp QL1 ( .CLK(CLK), .D(N_3), .PRE(CLR), .Q(ACO1) );

endmodule // upfxcar3

`endif

`ifdef upfxcar2
`else
`define upfxcar2
module upfxcar2( CLK , CLR, D, ENG, LOAD, ACO1, ACO2 );
output ACO1, ACO2;
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:1] D;
input ENG, LOAD;
supply0 GND;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
supply1 VCC;

mux4x7 QL8 ( .A(N_4), .B(N_4), .C(N_5), .D(ACO2), .Q(N_1), .S0(ENG), .S1(LOAD) );
mux4x7 QL7 ( .A(N_4), .B(N_4), .C(N_5), .D(ACO1), .Q(N_2), .S0(ENG), .S1(LOAD) );
upfxbit QL6 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENG(ENG), .ENP(GND), .ENT(GND),
           .LOAD(LOAD), .Q(N_3), .Q0(N_6), .Q1(VCC), .Q2(VCC) );
upfxbit QL5 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENG(ENG), .ENP(GND), .ENT(GND),
           .LOAD(LOAD), .Q(N_6), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
and2i1 QL4 ( .A(N_3), .B(N_6), .Q(N_5) );
and2i0 QL3 ( .A(D[0]), .B(D[1]), .Q(N_4) );
dffp QL2 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO2) );
dffp QL1 ( .CLK(CLK), .D(N_2), .PRE(CLR), .Q(ACO1) );

endmodule // upfxcar2

`endif

`ifdef upfxct4b
`else
`define upfxct4b
module upfxct4b( CLK , CLR, D, ENG, ENP, ENT, LOAD, Q, RCO );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:3] D;
input ENG, ENP, ENT, LOAD;
 output [0:3] Q;
output RCO;
supply1 VCC;

nand5i1 QL1 ( .A(Q[0]), .B(Q[1]), .C(Q[2]), .D(Q[3]), .E(ENT), .Q(RCO) );
upfxbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
upfxbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(VCC) );
upfxbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[1]), .Q0(Q[0]), .Q1(VCC), .Q2(VCC) );
upfxbit QL5 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[0]), .Q0(VCC), .Q1(VCC), .Q2(VCC) );

endmodule // upfxct4b

`endif

`ifdef upflcar1
`else
`define upflcar1
module upflcar1( CLK , CLR, D, LOAD, Q, ACO1 );
output ACO1;
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
 input [0:3] D;
input LOAD;
 input [0:3] Q;
supply0 GND;
supply1 VCC;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;

mux4x6 QL6 ( .A(VCC), .B(Q[3]), .C(D[3]), .D(VCC), .Q(N_1), .S0(N_4), .S1(N_5) );
and4i1 QL5 ( .A(LOAD), .B(N_3), .C(Q[2]), .D(N_2), .Q(N_4) );
and4i1 QL4 ( .A(D[0]), .B(D[1]), .C(D[2]), .D(LOAD), .Q(N_5) );
upflbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(N_3), .Q0(N_2), .Q1(VCC), .Q2(VCC) );
upflbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(N_2), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
dffp QL1 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO1) );

endmodule // upflcar1

`endif

`ifdef ucebit2a
`else
`define ucebit2a
module ucebit2a( CLK , CLR, ENH1, ENH2, ENH3, ENH4, ENL1, ENL2, ENL3, QFB, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input ENH1, ENH2, ENH3, ENH4, ENL1, ENL2, ENL3;
output Q;
input QFB;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

lcell2 I_1 ( .A1(ENH2), .A2(ENL3), .A3(ENH3), .A4(ENL2), .A5(ENH4), .A6(ENL1),
          .B1(GND), .B2(GND), .C1(QFB), .C2(GND), .D1(VCC), .D2(QFB), .E1(GND),
          .E2(GND), .F1(VCC), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND),
          .MP(GND), .MS(VCC), .NP(GND), .NS(GND), .OP(ENH1), .OS(GND), .QC(CLK),
          .QR(CLR), .QS(GND), .QZ(Q) );

endmodule // ucebit2a

`endif

`ifdef super_cell
`else
`define super_cell
module super_cell( A1 , A2, A3, A4, A5, A6, B1, B2, C1, C2, D1, D2, E1, E2, F1,
                   F2, F3, F4, F5, F6, MP, MS, NP, NS, OP, OS, PP, PS, QC, QR,
                   QS, AZ, FZ, NZ, OZ, Q2Z, QZ );
input A1, A2, A3, A4, A5, A6;
output AZ;
input B1, B2, C1, C2, D1, D2, E1, E2, F1, F2, F3, F4, F5, F6;
output FZ;
input MP, MS, NP, NS;
output NZ;
input OP, OS;
output OZ;
input PP, PS;
output Q2Z;
input QC;
input QR;
input QS;
output QZ;
parameter ql_frag = 1;
 wire TOPMUX_Z, MIDMUX_Z, BOTMUX_Z, FFMUX_Z, CLKMUX_Z; 
 wire MZ; 
 reg QZ, Q2Z; 
 
 assign #1 AZ = A1 & ~A2 & A3 & ~A4 & A5 & ~A6; 
 assign #1 TOPMUX_Z = OP ? AZ : OS; 
 assign #1 MZ = MIDMUX_Z ? (C1 & ~C2) : (B1 & ~B2); 
 assign #1 MIDMUX_Z = MP ? FZ : MS; 
 assign #1 NZ = BOTMUX_Z ? (E1 & ~E2) : (D1 & ~D2); 
 assign #1 BOTMUX_Z = NP ? FZ : NS; 
 assign #1 FZ = F1 & ~F2 & F3 & ~F4 & F5 & ~F6; 
 assign #1 OZ = TOPMUX_Z ? NZ : MZ; 
 assign #1 FFMUX_Z = PP ? PS : NZ; 
`ifdef synthesis 
  always @ (posedge QC or posedge QR or posedge QS) 
     if (QR) 
        #1 QZ = 1'b0; 
     else if (QS) 
        #1 QZ = 1'b1; 
     else 
        #1 QZ = OZ; 
  always @ (posedge QC or posedge QR or posedge QS) 
     if (QR) 
        #1 Q2Z = 1'b0; 
     else if (QS) 
        #1 Q2Z = 1'b1; 
     else 
        #1 Q2Z = FFMUX_Z; 
`else 
  always @ (posedge QC) 
     if (~QR && ~QS) 
        #1 QZ = OZ; 
  always @ (QR or QS) 
     if (QR) 
        #1 QZ = 1'b0; 
     else if (QS) 
        #1 QZ = 1'b1; 
  always @ (posedge QC) 
     if (~QR && ~QS) 
        #1 Q2Z = FFMUX_Z; 
  always @ (QR or QS) 
     if (QR) 
        #1 Q2Z = 1'b0; 
     else if (QS) 
        #1 Q2Z = 1'b1; 
`endif 

endmodule // super_cell

`endif

`ifdef hsckmux
`else
`define hsckmux
module hsckmux( IC , IS, IZ );
input IC, IS;
output IZ;
parameter ql_frag = 1;
 assign #1 IZ = IS ? IC : 1'b0;

endmodule // hsckmux

`endif

`ifdef eio_cell
`else
`define eio_cell
module eio_cell( EQE , ESEL, IE, IQC, IQE, IQR, OQI, OSEL, IQQ, IZ, OQQ, IP );
input EQE;
input ESEL, IE;
inout IP;
input IQC;
input IQE;
output IQQ;
input IQR;
output IZ;
input OQI;
output OQQ;
input OSEL;
parameter ql_frag = 1;
 wire EQMUX_Z, OQMUX_Z; 
 reg EQZ, OQQ, IQQ; 
 assign #1 EQMUX_Z = ESEL ? IE : EQZ; 
 assign #1 OQMUX_Z = OSEL ? OQI : OQQ; 
 assign #1 IP = EQMUX_Z ? OQMUX_Z : 1'bz; 
 assign #1 IZ = IP; 
`ifdef synthesis 
  always @ (posedge IQC or posedge IQR) 
    if (IQR)
      #1 EQZ = 1'b0;
    else if (EQE)
      #1 EQZ = IE; 
  always @ (posedge IQC or posedge IQR) 
    if (IQR)
      #1 IQQ = 1'b0; 
    else if (IQE) 
      #1 IQQ = IP; 
  always @ (posedge IQC or posedge IQR) 
    if (IQR) 
      #1 OQQ = 1'b0; 
    else 
      #1 OQQ = OQI; 
`else 
  always @ (posedge IQC) 
    if (~IQR & EQE)
      #1 EQZ = IE; 
    else if (IQR) 
      #1 EQZ = 1'b0;
  always @ (posedge IQC) 
    if (~IQR & IQE) 
      #1 IQQ = IP; 
    else if (IQR) 
      #1 IQQ = 1'b0;  always @ (posedge IQC) 
    if (~IQR) 
      #1 OQQ = OQI; 
    else if (IQR) 
      #1 OQQ = 1'b0; 
`endif 

endmodule // eio_cell

`endif

`ifdef inbuffcell_25um
`else
`define inbuffcell_25um
module inbuffcell_25um( I, IP, IS, O );
input I, IP, IS;
output O;
parameter ql_frag = 1;
 assign #1 O = IS ? I : IP; 

endmodule // inbuffcell_25um

`endif

`ifdef iocontrol
`else
`define iocontrol
module iocontrol( IP , IS, O );
input IP, IS;
output O;
parameter ql_frag = 1;
 assign #1 O = IS ? 1'b0 : IP; 

endmodule // iocontrol

`endif

`ifdef ckcell_25um
`else
`define ckcell_25um
module ckcell_25um( IP , IC );
output IC;
input IP;
parameter ql_frag = 1;
 assign #1 IC = IP;

endmodule // ckcell_25um

`endif

`ifdef ckcell5
`else
`define ckcell5
module ckcell5( IP , IC );
output IC;
input IP;
parameter ql_frag = 1;
 assign #1 IC = IP;

endmodule // ckcell5

`endif

`ifdef lcell2
`else
`define lcell2
module lcell2( A1 , A2, A3, A4, A5, A6, B1, B2, C1, C2, D1, D2, E1, E2, F1, F2,
               F3, F4, F5, F6, MP, MS, NP, NS, OP, OS, QC, QR, QS, AZ, FZ, NZ,
               OZ, QZ );
input A1, A2, A3, A4, A5, A6;
output AZ;
input B1, B2, C1, C2, D1, D2, E1, E2, F1, F2, F3, F4, F5, F6;
output FZ;
input MP, MS, NP, NS;
output NZ;
input OP, OS;
output OZ;
input QC, QR, QS;
output QZ;
parameter syn_macro = 1, ql_pack = 1;
parameter ql_frag = 1;
 wire TOPMUX_Z, MIDMUX_Z, BOTMUX_Z; 
 wire MZ; 
 reg QZ; 
 
 assign #1 AZ = A1 & ~A2 & A3 & ~A4 & A5 & ~A6; 
 assign #1 TOPMUX_Z = OP ? AZ : OS;  
 assign #1 MZ = MIDMUX_Z ? (C1 & ~C2):(B1 & ~B2); 
 assign #1 MIDMUX_Z = MP ? FZ : MS;  
 assign #1 NZ = BOTMUX_Z ? (E1 & ~E2):(D1 & ~D2); 
 assign #1 BOTMUX_Z = NP ? FZ : NS;  
 assign #1 FZ = F1 & ~F2 & F3 & ~F4 & F5 & ~F6; 
 assign #1 OZ = TOPMUX_Z ? NZ : MZ;  
`ifdef synthesis 
 always @ (posedge QC or posedge QR or posedge QS)  
     if (QR) 
        #1 QZ = 1'b0; 
     else if (QS) 
        #1 QZ = 1'b1; 
     else #1 QZ = OZ; 
`else 
  always @ (posedge QC) 
      if (~QR && ~QS) 
         #1 QZ = OZ; 
  always @ (QR or QS) 
      if (QR) 
         #1 QZ = 1'b0; 
      else if (QS) 
         #1 QZ = 1'b1; 
 `endif 

endmodule // lcell2

`endif

`ifdef ucxco
`else
`define ucxco
module ucxco( CLK , D_DEC, EN, LOAD, PRE, Q_DEC, CO, LDBUF );
input CLK /* synthesis syn_isclock=1 */;
output CO;
input D_DEC, EN;
output LDBUF;
input PRE /* synthesis syn_isclock=1 */;
input LOAD, Q_DEC;
parameter ql_gate = `LOGIC;
supply0 GND;
supply1 VCC;

lcell2 I_1 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(LOAD),
          .AZ(LDBUF), .B1(VCC), .B2(Q_DEC), .C1(CO), .C2(GND), .D1(VCC),
          .D2(D_DEC), .E1(GND), .E2(GND), .F1(VCC), .F2(GND), .F3(VCC), .F4(GND),
          .F5(VCC), .F6(GND), .MP(GND), .MS(EN), .NP(GND), .NS(GND), .OP(VCC),
          .OS(GND), .QC(CLK), .QR(GND), .QS(PRE), .QZ(CO) );

endmodule // ucxco

`endif

`ifdef ucxbit2b
`else
`define ucxbit2b
module ucxbit2b( CLK , CLR, D, ENH1, ENH2, ENH3, ENH4, ENL1, ENL2, ENL3, LOAD,
                 QFB, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input D, ENH1, ENH2, ENH3, ENH4, ENL1, ENL2, ENL3, LOAD;
output Q;
input QFB;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

lcell2 I_2 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .B1(VCC),
          .B2(QFB), .C1(QFB), .C2(GND), .D1(D), .D2(GND), .E1(GND), .E2(GND),
          .F1(ENH2), .F2(ENL3), .F3(ENH3), .F4(ENL2), .F5(ENH4), .F6(ENL1),
          .MP(ENH1), .MS(GND), .NP(GND), .NS(GND), .OP(GND), .OS(LOAD), .QC(CLK),
          .QR(CLR), .QS(GND), .QZ(Q) );

endmodule // ucxbit2b

`endif

`ifdef ucxbit2a
`else
`define ucxbit2a
module ucxbit2a( CLK , CLR, D, ENH1, ENH2, ENH3, ENH4, ENL1, ENL2, ENL3, LOAD,
                 QFB, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input D, ENH1, ENH2, ENH3, ENH4, ENL1, ENL2, ENL3, LOAD;
output Q;
input QFB;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

lcell2 I_2 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .B1(QFB),
          .B2(GND), .C1(VCC), .C2(QFB), .D1(D), .D2(GND), .E1(GND), .E2(GND),
          .F1(ENH2), .F2(ENL3), .F3(ENH3), .F4(ENL2), .F5(ENH4), .F6(ENL1),
          .MP(ENH1), .MS(GND), .NP(GND), .NS(GND), .OP(GND), .OS(LOAD), .QC(CLK),
          .QR(CLR), .QS(GND), .QZ(Q) );

endmodule // ucxbit2a

`endif

`ifdef dif32
`else
`define dif32
module dif32( a , b, C11_C70, C11_C71, C19_C150, C19_C151, C23_C190, C23_C191,
              C27_C230, C27_C231, C7_C30, C7_C31, Carry15, Carry15a, Carry15b,
              Cin, Co0_Ci0, Co0_Ci1, Co10_C90, Co10_C91, Co12_C110, Co12_C111,
              Co13_C120, Co13_C121, Co14_C130, Co14_C131, Co16_C150,
              Co16_C151, Co17_C160, Co17_C161, Co18_C170, Co18_C171, Co1_C00,
              Co1_C01, Co20_C190, Co20_C191, Co21_C200, Co21_C201, Co22_C210,
              Co22_C211, Co24_C230, Co24_C231, Co25_C240, Co25_C241,
              Co26_C250, Co26_C251, Co28_C270, Co28_C271, Co29_C280,
              Co29_C281, Co2_C10, Co2_C11, Co30_C290, Co30_C291, Co3_C20,
              Co3_C21, Co4_C30, Co4_C31, Co5_C40, Co5_C41, Co6_C50, Co6_C51,
              Co8_C70, Co8_C71, Co9_C80, Co9_C81, S, Carry3, Carry3a, Sumi );
 input [0:0] a;
 input [0:0] b;
input C11_C70, C11_C71, C19_C150, C19_C151, C23_C190, C23_C191, C27_C230,
C27_C231, C7_C30, C7_C31, Carry15, Carry15a, Carry15b;
output Carry3, Carry3a;
input Cin, Co0_Ci0, Co0_Ci1, Co10_C90, Co10_C91, Co12_C110, Co12_C111,
Co13_C120, Co13_C121, Co14_C130, Co14_C131, Co16_C150, Co16_C151,
Co17_C160, Co17_C161, Co18_C170, Co18_C171, Co1_C00, Co1_C01,
Co20_C190, Co20_C191, Co21_C200, Co21_C201, Co22_C210, Co22_C211,
Co24_C230, Co24_C231, Co25_C240, Co25_C241, Co26_C250, Co26_C251,
Co28_C270, Co28_C271, Co29_C280, Co29_C281, Co2_C10, Co2_C11,
Co30_C290, Co30_C291, Co3_C20, Co3_C21, Co4_C30, Co4_C31, Co5_C40,
Co5_C41, Co6_C50, Co6_C51, Co8_C70, Co8_C71, Co9_C80, Co9_C81;
 input [31:0] S;
 output [31:0] Sumi;
wire N_189;
wire N_190;
wire N_191;
wire N_192;
wire N_193;
wire N_194;
wire N_195;
wire N_196;
wire N_197;
wire N_198;
wire N_199;
wire N_200;
wire N_181;
wire N_182;
wire N_183;
wire N_184;
wire N_185;
wire N_186;
wire N_187;
wire N_188;
wire N_175;
wire N_180;
wire N_135;
wire N_139;
wire N_152;
wire N_153;
wire N_94;
wire N_95;
wire N_41;
wire N_42;
wire N_43;
wire N_44;
wire N_40;
wire N_37;
wire Carry0;
supply0 gnd;

borrow0 I_135 ( .A(a[0]), .B(b[0]), .Bin(Cin), .Bout(Carry0) );
dif0 I_134 ( .A(a[0]), .B(b[0]), .Bin(Cin), .d0(Sumi[0]) );
mux2x0 I_133 ( .A(N_187), .B(N_188), .Q(Sumi[31]), .S(Carry15b) );
sum2_gen I161 ( .C_i(C19_C151), .Cj_i0(C23_C190), .Cj_i1(C23_C191),
             .Ck_j0(C27_C230), .Ck_j1(C27_C231), .Sk_0(N_185), .Sk_1(N_186),
             .Sk_i(N_188) );
sum2_gen I_122 ( .C_i(C19_C150), .Cj_i0(C23_C190), .Cj_i1(C23_C191),
              .Ck_j0(C27_C230), .Ck_j1(C27_C231), .Sk_0(N_185), .Sk_1(N_186),
              .Sk_i(N_187) );
sum2_gen I_129 ( .C_i(Carry15b), .Cj_i0(C19_C150), .Cj_i1(C19_C151),
              .Ck_j0(C23_C190), .Ck_j1(C23_C191), .Sk_0(N_139), .Sk_1(N_135),
              .Sk_i(Sumi[30]) );
sum2_gen I162 ( .C_i(Carry15b), .Cj_i0(C19_C150), .Cj_i1(C19_C151),
             .Ck_j0(C23_C190), .Ck_j1(C23_C191), .Sk_0(N_153), .Sk_1(N_152),
             .Sk_i(Sumi[29]) );
sum2_gen I_119 ( .C_i(Carry15a), .Cj_i0(C19_C150), .Cj_i1(C19_C151),
              .Ck_j0(C23_C190), .Ck_j1(C23_C191), .Sk_0(N_94), .Sk_1(N_95),
              .Sk_i(Sumi[28]) );
sum2_gen I_106 ( .C_i(Carry15b), .Cj_i0(C19_C150), .Cj_i1(C19_C151),
              .Ck_j0(C23_C190), .Ck_j1(C23_C191), .Sk_0(N_40), .Sk_1(N_37),
              .Sk_i(Sumi[25]) );
sum2_gen I_107 ( .C_i(Carry15b), .Cj_i0(C19_C150), .Cj_i1(C19_C151),
              .Ck_j0(C23_C190), .Ck_j1(C23_C191), .Sk_0(N_44), .Sk_1(N_43),
              .Sk_i(Sumi[26]) );
sum2_gen I_108 ( .C_i(Carry15b), .Cj_i0(C19_C150), .Cj_i1(C19_C151),
              .Ck_j0(C23_C190), .Ck_j1(C23_C191), .Sk_0(N_42), .Sk_1(N_41),
              .Sk_i(Sumi[27]) );
sum2_gen I_99 ( .C_i(gnd), .Cj_i0(Carry15), .Cj_i1(gnd), .Ck_j0(C19_C150),
             .Ck_j1(C19_C151), .Sk_0(N_184), .Sk_1(N_182), .Sk_i(Sumi[23]) );
sum2_gen I_100 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Carry15),
              .Ck_j1(gnd), .Sk_0(N_183), .Sk_1(N_181), .Sk_i(Sumi[22]) );
sum2_gen I_90 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Carry15a),
             .Ck_j1(gnd), .Sk_0(N_180), .Sk_1(N_175), .Sk_i(Sumi[19]) );
sum2_gen I153 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Carry3), .Ck_j1(gnd),
             .Sk_0(N_189), .Sk_1(N_190), .Sk_i(Sumi[7]) );
sum2_gen I154 ( .C_i(Carry3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
             .Ck_j1(C11_C71), .Sk_0(N_200), .Sk_1(N_197), .Sk_i(Sumi[15]) );
sum2_gen I155 ( .C_i(Carry3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
             .Ck_j1(C11_C71), .Sk_0(N_198), .Sk_1(N_196), .Sk_i(Sumi[14]) );
sum2_gen I156 ( .C_i(Carry3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
             .Ck_j1(C11_C71), .Sk_0(N_199), .Sk_1(N_195), .Sk_i(Sumi[13]) );
sum2_gen I157 ( .C_i(gnd), .Cj_i0(Carry3a), .Cj_i1(gnd), .Ck_j0(C7_C30),
             .Ck_j1(C7_C31), .Sk_0(N_194), .Sk_1(N_191), .Sk_i(Sumi[11]) );
sum2_gen I158 ( .C_i(gnd), .Cj_i0(Carry3a), .Cj_i1(gnd), .Ck_j0(C7_C30),
             .Ck_j1(C7_C31), .Sk_0(N_192), .Sk_1(N_193), .Sk_i(Sumi[10]) );
cary_gen I159 ( .C_i(Carry0), .Cj_i0(Co1_C00), .Cj_i1(Co1_C01), .Ck_j0(Co2_C10),
             .Ck_j1(Co2_C11), .Cm_i(Carry3a), .Cm_k0(Co3_C20),
             .Cm_k1(Co3_C21) );
cary_gen I160 ( .C_i(Carry0), .Cj_i0(Co1_C00), .Cj_i1(Co1_C01), .Ck_j0(Co2_C10),
             .Ck_j1(Co2_C11), .Cm_i(Carry3), .Cm_k0(Co3_C20), .Cm_k1(Co3_C21) );
sum_gen I163 ( .C_i(Co28_C271), .Cj_i0(Co29_C280), .Cj_i1(Co29_C281),
            .Ck_j0(Co30_C290), .Ck_j1(Co30_C291), .Sk_01(S[31]), .Sk_i(N_186) );
sum_gen I_125 ( .C_i(Co28_C270), .Cj_i0(Co29_C280), .Cj_i1(Co29_C281),
             .Ck_j0(Co30_C290), .Ck_j1(Co30_C291), .Sk_01(S[31]),
             .Sk_i(N_185) );
sum_gen I164 ( .C_i(C27_C231), .Cj_i0(Co28_C270), .Cj_i1(Co28_C271),
            .Ck_j0(Co29_C280), .Ck_j1(Co29_C281), .Sk_01(S[30]), .Sk_i(N_135) );
sum_gen I_131 ( .C_i(C27_C230), .Cj_i0(Co28_C270), .Cj_i1(Co28_C271),
             .Ck_j0(Co29_C280), .Ck_j1(Co29_C281), .Sk_01(S[30]),
             .Sk_i(N_139) );
sum_gen I165 ( .C_i(gnd), .Cj_i0(C27_C231), .Cj_i1(gnd), .Ck_j0(Co28_C270),
            .Ck_j1(Co28_C271), .Sk_01(S[29]), .Sk_i(N_152) );
sum_gen I166 ( .C_i(gnd), .Cj_i0(C27_C230), .Cj_i1(gnd), .Ck_j0(Co28_C270),
            .Ck_j1(Co28_C271), .Sk_01(S[29]), .Sk_i(N_153) );
sum_gen I167 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(C27_C231), .Ck_j1(gnd),
            .Sk_01(S[28]), .Sk_i(N_95) );
sum_gen I_120 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(C27_C230),
             .Ck_j1(gnd), .Sk_01(S[28]), .Sk_i(N_94) );
sum_gen I168 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Co24_C231),
            .Ck_j1(gnd), .Sk_01(S[25]), .Sk_i(N_37) );
sum_gen I169 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Co24_C230),
            .Ck_j1(gnd), .Sk_01(S[25]), .Sk_i(N_40) );
sum_gen I_105 ( .C_i(Carry15), .Cj_i0(C19_C150), .Cj_i1(C19_C151),
             .Ck_j0(C23_C190), .Ck_j1(C23_C191), .Sk_01(S[24]),
             .Sk_i(Sumi[24]) );
sum_gen I_102 ( .C_i(gnd), .Cj_i0(Co24_C230), .Cj_i1(gnd), .Ck_j0(Co25_C240),
             .Ck_j1(Co25_C241), .Sk_01(S[26]), .Sk_i(N_44) );
sum_gen I170 ( .C_i(Co24_C231), .Cj_i0(Co25_C240), .Cj_i1(Co25_C241),
            .Ck_j0(Co26_C250), .Ck_j1(Co26_C251), .Sk_01(S[27]), .Sk_i(N_41) );
sum_gen I171 ( .C_i(Co24_C230), .Cj_i0(Co25_C240), .Cj_i1(Co25_C241),
            .Ck_j0(Co26_C250), .Ck_j1(Co26_C251), .Sk_01(S[27]), .Sk_i(N_42) );
sum_gen I_101 ( .C_i(gnd), .Cj_i0(Co24_C231), .Cj_i1(gnd), .Ck_j0(Co25_C240),
             .Ck_j1(Co25_C241), .Sk_01(S[26]), .Sk_i(N_43) );
sum_gen I_93 ( .C_i(Co20_C191), .Cj_i0(Co21_C200), .Cj_i1(Co21_C201),
            .Ck_j0(Co22_C210), .Ck_j1(Co22_C211), .Sk_01(S[23]), .Sk_i(N_182) );
sum_gen I_92 ( .C_i(Co20_C190), .Cj_i0(Co21_C200), .Cj_i1(Co21_C201),
            .Ck_j0(Co22_C210), .Ck_j1(Co22_C211), .Sk_01(S[23]), .Sk_i(N_184) );
sum_gen I_94 ( .C_i(C19_C151), .Cj_i0(Co20_C190), .Cj_i1(Co20_C191),
            .Ck_j0(Co21_C200), .Ck_j1(Co21_C201), .Sk_01(S[22]), .Sk_i(N_181) );
sum_gen I_95 ( .C_i(C19_C150), .Cj_i0(Co20_C190), .Cj_i1(Co20_C191),
            .Ck_j0(Co21_C200), .Ck_j1(Co21_C201), .Sk_01(S[22]), .Sk_i(N_183) );
sum_gen I_91 ( .C_i(Carry15), .Cj_i0(C19_C150), .Cj_i1(C19_C151),
            .Ck_j0(Co20_C190), .Ck_j1(Co20_C191), .Sk_01(S[21]),
            .Sk_i(Sumi[21]) );
sum_gen I_97 ( .C_i(gnd), .Cj_i0(Carry15), .Cj_i1(gnd), .Ck_j0(C19_C150),
            .Ck_j1(C19_C151), .Sk_01(S[20]), .Sk_i(Sumi[20]) );
sum_gen I_89 ( .C_i(Co16_C151), .Cj_i0(Co17_C160), .Cj_i1(Co17_C161),
            .Ck_j0(Co18_C170), .Ck_j1(Co18_C171), .Sk_01(S[19]), .Sk_i(N_175) );
sum_gen I_84 ( .C_i(Co16_C150), .Cj_i0(Co17_C160), .Cj_i1(Co17_C161),
            .Ck_j0(Co18_C170), .Ck_j1(Co18_C171), .Sk_01(S[19]), .Sk_i(N_180) );
sum_gen I_85 ( .C_i(Carry15a), .Cj_i0(Co16_C150), .Cj_i1(Co16_C151),
            .Ck_j0(Co17_C160), .Ck_j1(Co17_C161), .Sk_01(S[18]),
            .Sk_i(Sumi[18]) );
sum_gen I_86 ( .C_i(gnd), .Cj_i0(Carry15a), .Cj_i1(gnd), .Ck_j0(Co16_C150),
            .Ck_j1(Co16_C151), .Sk_01(S[17]), .Sk_i(Sumi[17]) );
sum_gen I_87 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Carry15a), .Ck_j1(gnd),
            .Sk_01(S[16]), .Sk_i(Sumi[16]) );
sum_gen sum15_1 ( .C_i(Co12_C111), .Cj_i0(Co13_C120), .Cj_i1(Co13_C121),
               .Ck_j0(Co14_C130), .Ck_j1(Co14_C131), .Sk_01(S[15]),
               .Sk_i(N_197) );
sum_gen I147 ( .C_i(Co12_C110), .Cj_i0(Co13_C120), .Cj_i1(Co13_C121),
            .Ck_j0(Co14_C130), .Ck_j1(Co14_C131), .Sk_01(S[15]), .Sk_i(N_200) );
sum_gen I148 ( .C_i(gnd), .Cj_i0(Co12_C111), .Cj_i1(gnd), .Ck_j0(Co13_C120),
            .Ck_j1(Co13_C121), .Sk_01(S[14]), .Sk_i(N_196) );
sum_gen I149 ( .C_i(gnd), .Cj_i0(Co12_C110), .Cj_i1(gnd), .Ck_j0(Co13_C120),
            .Ck_j1(Co13_C121), .Sk_01(S[14]), .Sk_i(N_198) );
sum_gen I150 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Co12_C111),
            .Ck_j1(gnd), .Sk_01(S[13]), .Sk_i(N_195) );
sum_gen I151 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Co12_C110),
            .Ck_j1(gnd), .Sk_01(S[13]), .Sk_i(N_199) );
sum_gen I152 ( .C_i(Carry3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
            .Ck_j1(C11_C71), .Sk_01(S[12]), .Sk_i(Sumi[12]) );
sum_gen I133 ( .C_i(Co4_C31), .Cj_i0(Co5_C40), .Cj_i1(Co5_C41), .Ck_j0(Co6_C50),
            .Ck_j1(Co6_C51), .Sk_01(S[7]), .Sk_i(N_190) );
sum_gen I134 ( .C_i(Co4_C30), .Cj_i0(Co5_C40), .Cj_i1(Co5_C41), .Ck_j0(Co6_C50),
            .Ck_j1(Co6_C51), .Sk_01(S[7]), .Sk_i(N_189) );
sum_gen I135 ( .C_i(Carry3), .Cj_i0(Co4_C30), .Cj_i1(Co4_C31), .Ck_j0(Co5_C40),
            .Ck_j1(Co5_C41), .Sk_01(S[6]), .Sk_i(Sumi[6]) );
sum_gen I136 ( .C_i(gnd), .Cj_i0(Carry3), .Cj_i1(gnd), .Ck_j0(Co4_C30),
            .Ck_j1(Co4_C31), .Sk_01(S[5]), .Sk_i(Sumi[5]) );
sum_gen I137 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Carry3), .Ck_j1(gnd),
            .Sk_01(S[4]), .Sk_i(Sumi[4]) );
sum_gen I138 ( .C_i(Co8_C71), .Cj_i0(Co9_C80), .Cj_i1(Co9_C81), .Ck_j0(Co10_C90),
            .Ck_j1(Co10_C91), .Sk_01(S[11]), .Sk_i(N_191) );
sum_gen I139 ( .C_i(Co8_C70), .Cj_i0(Co9_C80), .Cj_i1(Co9_C81), .Ck_j0(Co10_C90),
            .Ck_j1(Co10_C91), .Sk_01(S[11]), .Sk_i(N_194) );
sum_gen I140 ( .C_i(gnd), .Cj_i0(Co8_C71), .Cj_i1(gnd), .Ck_j0(Co9_C80),
            .Ck_j1(Co9_C81), .Sk_01(S[10]), .Sk_i(N_193) );
sum_gen I141 ( .C_i(gnd), .Cj_i0(Co8_C70), .Cj_i1(gnd), .Ck_j0(Co9_C80),
            .Ck_j1(Co9_C81), .Sk_01(S[10]), .Sk_i(N_192) );
sum_gen I142 ( .C_i(Carry3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(Co8_C70),
            .Ck_j1(Co8_C71), .Sk_01(S[9]), .Sk_i(Sumi[9]) );
sum_gen I143 ( .C_i(gnd), .Cj_i0(Carry3a), .Cj_i1(gnd), .Ck_j0(C7_C30),
            .Ck_j1(C7_C31), .Sk_01(S[8]), .Sk_i(Sumi[8]) );
sum_gen I144 ( .C_i(Carry0), .Cj_i0(Co1_C00), .Cj_i1(Co1_C01), .Ck_j0(Co2_C10),
            .Ck_j1(Co2_C11), .Sk_01(S[3]), .Sk_i(Sumi[3]) );
sum_gen I145 ( .C_i(Cin), .Cj_i0(Co0_Ci1), .Cj_i1(Co0_Ci0), .Ck_j0(Co1_C00),
            .Ck_j1(Co1_C01), .Sk_01(S[2]), .Sk_i(Sumi[2]) );
sum_gen I146 ( .C_i(gnd), .Cj_i0(Cin), .Cj_i1(gnd), .Ck_j0(Co0_Ci1),
            .Ck_j1(Co0_Ci0), .Sk_01(S[1]), .Sk_i(Sumi[1]) );

endmodule // dif32

`endif

`ifdef borrow32
`else
`define borrow32
module borrow32( a , b, Carry3, Carry3a, C11_C70, C11_C71, C19_C150, C19_C151,
                 C23_C190, C23_C191, C27_C230, C27_C231, C7_C30, C7_C31,
                 Carry15, Carry15a, Carry15b, Co, Co0_Ci0, Co0_Ci1, Co10_C90,
                 Co10_C91, Co12_C110, Co12_C111, Co13_C120, Co13_C121,
                 Co14_C130, Co14_C131, Co16_C150, Co16_C151, Co17_C160,
                 Co17_C161, Co18_C170, Co18_C171, Co1_C00, Co1_C01, Co20_C190,
                 Co20_C191, Co21_C200, Co21_C201, Co22_C210, Co22_C211,
                 Co24_C230, Co24_C231, Co25_C240, Co25_C241, Co26_C250,
                 Co26_C251, Co28_C270, Co28_C271, Co29_C280, Co29_C281,
                 Co2_C10, Co2_C11, Co30_C290, Co30_C291, Co3_C20, Co3_C21,
                 Co4_C30, Co4_C31, Co5_C40, Co5_C41, Co6_C50, Co6_C51,
                 Co8_C70, Co8_C71, Co9_C80, Co9_C81, S );
 input [31:0] a;
 input [31:0] b;
output C11_C70, C11_C71, C19_C150, C19_C151, C23_C190, C23_C191, C27_C230,
C27_C231, C7_C30, C7_C31, Carry15, Carry15a, Carry15b;
input Carry3, Carry3a;
output Co, Co0_Ci0, Co0_Ci1, Co10_C90, Co10_C91, Co12_C110, Co12_C111,
Co13_C120, Co13_C121, Co14_C130, Co14_C131, Co16_C150, Co16_C151,
Co17_C160, Co17_C161, Co18_C170, Co18_C171, Co1_C00, Co1_C01,
Co20_C190, Co20_C191, Co21_C200, Co21_C201, Co22_C210, Co22_C211,
Co24_C230, Co24_C231, Co25_C240, Co25_C241, Co26_C250, Co26_C251,
Co28_C270, Co28_C271, Co29_C280, Co29_C281, Co2_C10, Co2_C11,
Co30_C290, Co30_C291, Co3_C20, Co3_C21, Co4_C30, Co4_C31, Co5_C40,
Co5_C41, Co6_C50, Co6_C51, Co8_C70, Co8_C71, Co9_C80, Co9_C81;
 output [31:0] S;
wire C31_C160;
wire C31_C161;
wire Co19_C180;
wire Co19_C181;
wire Co23_C220;
wire Co23_C221;
wire Co27_C260;
wire Co27_C261;
wire Co31_C300;
wire Co31_C301;
wire Co7_C60;
wire Co7_C61;
wire Co11_C100;
wire Co11_C101;
wire Co15_C140;
wire Co15_C141;
wire C31_C270;
wire C31_C271;
wire C15_C110;
wire C15_C111;

dif_b0 I_106 ( .Ax(a[0]), .Bo_Bi0(Co0_Ci0), .Bo_Bi1(Co0_Ci1), .Bx(b[0]) );
dif_b I_89 ( .Ax(a[16]), .Bo_Bi0(Co16_C150), .Bo_Bi1(Co16_C151), .Bx(b[16]),
          .Sub_Dif(S[16]) );
dif_b I_88 ( .Ax(a[17]), .Bo_Bi0(Co17_C160), .Bo_Bi1(Co17_C161), .Bx(b[17]),
          .Sub_Dif(S[17]) );
dif_b I_87 ( .Ax(a[18]), .Bo_Bi0(Co18_C170), .Bo_Bi1(Co18_C171), .Bx(b[18]),
          .Sub_Dif(S[18]) );
dif_b I_86 ( .Ax(a[19]), .Bo_Bi0(Co19_C180), .Bo_Bi1(Co19_C181), .Bx(b[19]),
          .Sub_Dif(S[19]) );
dif_b I_85 ( .Ax(a[20]), .Bo_Bi0(Co20_C190), .Bo_Bi1(Co20_C191), .Bx(b[20]),
          .Sub_Dif(S[20]) );
dif_b I_84 ( .Ax(a[21]), .Bo_Bi0(Co21_C200), .Bo_Bi1(Co21_C201), .Bx(b[21]),
          .Sub_Dif(S[21]) );
dif_b I_83 ( .Ax(a[22]), .Bo_Bi0(Co22_C210), .Bo_Bi1(Co22_C211), .Bx(b[22]),
          .Sub_Dif(S[22]) );
dif_b I_82 ( .Ax(a[23]), .Bo_Bi0(Co23_C220), .Bo_Bi1(Co23_C221), .Bx(b[23]),
          .Sub_Dif(S[23]) );
dif_b I_81 ( .Ax(a[24]), .Bo_Bi0(Co24_C230), .Bo_Bi1(Co24_C231), .Bx(b[24]),
          .Sub_Dif(S[24]) );
dif_b I_80 ( .Ax(a[25]), .Bo_Bi0(Co25_C240), .Bo_Bi1(Co25_C241), .Bx(b[25]),
          .Sub_Dif(S[25]) );
dif_b I_79 ( .Ax(a[26]), .Bo_Bi0(Co26_C250), .Bo_Bi1(Co26_C251), .Bx(b[26]),
          .Sub_Dif(S[26]) );
dif_b I_78 ( .Ax(a[27]), .Bo_Bi0(Co27_C260), .Bo_Bi1(Co27_C261), .Bx(b[27]),
          .Sub_Dif(S[27]) );
dif_b I_77 ( .Ax(a[28]), .Bo_Bi0(Co28_C270), .Bo_Bi1(Co28_C271), .Bx(b[28]),
          .Sub_Dif(S[28]) );
dif_b I_76 ( .Ax(a[29]), .Bo_Bi0(Co29_C280), .Bo_Bi1(Co29_C281), .Bx(b[29]),
          .Sub_Dif(S[29]) );
dif_b I_75 ( .Ax(a[30]), .Bo_Bi0(Co30_C290), .Bo_Bi1(Co30_C291), .Bx(b[30]),
          .Sub_Dif(S[30]) );
dif_b I_74 ( .Ax(a[31]), .Bo_Bi0(Co31_C300), .Bo_Bi1(Co31_C301), .Bx(b[31]),
          .Sub_Dif(S[31]) );
dif_b I_105 ( .Ax(a[1]), .Bo_Bi0(Co1_C00), .Bo_Bi1(Co1_C01), .Bx(b[1]),
           .Sub_Dif(S[1]) );
dif_b I_103 ( .Ax(a[2]), .Bo_Bi0(Co2_C10), .Bo_Bi1(Co2_C11), .Bx(b[2]),
           .Sub_Dif(S[2]) );
dif_b I_102 ( .Ax(a[3]), .Bo_Bi0(Co3_C20), .Bo_Bi1(Co3_C21), .Bx(b[3]),
           .Sub_Dif(S[3]) );
dif_b I_101 ( .Ax(a[4]), .Bo_Bi0(Co4_C30), .Bo_Bi1(Co4_C31), .Bx(b[4]),
           .Sub_Dif(S[4]) );
dif_b I_100 ( .Ax(a[5]), .Bo_Bi0(Co5_C40), .Bo_Bi1(Co5_C41), .Bx(b[5]),
           .Sub_Dif(S[5]) );
dif_b I_99 ( .Ax(a[6]), .Bo_Bi0(Co6_C50), .Bo_Bi1(Co6_C51), .Bx(b[6]),
          .Sub_Dif(S[6]) );
dif_b I_98 ( .Ax(a[7]), .Bo_Bi0(Co7_C60), .Bo_Bi1(Co7_C61), .Bx(b[7]),
          .Sub_Dif(S[7]) );
dif_b I_97 ( .Ax(a[8]), .Bo_Bi0(Co8_C70), .Bo_Bi1(Co8_C71), .Bx(b[8]),
          .Sub_Dif(S[8]) );
dif_b I_96 ( .Ax(a[9]), .Bo_Bi0(Co9_C80), .Bo_Bi1(Co9_C81), .Bx(b[9]),
          .Sub_Dif(S[9]) );
dif_b I_95 ( .Ax(a[10]), .Bo_Bi0(Co10_C90), .Bo_Bi1(Co10_C91), .Bx(b[10]),
          .Sub_Dif(S[10]) );
dif_b I_94 ( .Ax(a[11]), .Bo_Bi0(Co11_C100), .Bo_Bi1(Co11_C101), .Bx(b[11]),
          .Sub_Dif(S[11]) );
dif_b I_93 ( .Ax(a[12]), .Bo_Bi0(Co12_C110), .Bo_Bi1(Co12_C111), .Bx(b[12]),
          .Sub_Dif(S[12]) );
dif_b I_91 ( .Ax(a[14]), .Bo_Bi0(Co14_C130), .Bo_Bi1(Co14_C131), .Bx(b[14]),
          .Sub_Dif(S[14]) );
dif_b I_90 ( .Ax(a[15]), .Bo_Bi0(Co15_C140), .Bo_Bi1(Co15_C141), .Bx(b[15]),
          .Sub_Dif(S[15]) );
dif_b I_92 ( .Ax(a[13]), .Bo_Bi0(Co13_C120), .Bo_Bi1(Co13_C121), .Bx(b[13]),
          .Sub_Dif(S[13]) );
b_out I_73 ( .Bo(Co), .By_x0(Carry15), .Bz_y0(C31_C160), .Bz_y1(C31_C161) );
cary_gen I104 ( .C_i(Co12_C111), .Cj_i0(Co13_C120), .Cj_i1(Co13_C121),
             .Ck_j0(Co14_C130), .Ck_j1(Co14_C131), .Cm_i(C15_C111),
             .Cm_k0(Co15_C140), .Cm_k1(Co15_C141) );
cary_gen I105 ( .C_i(Co12_C110), .Cj_i0(Co13_C120), .Cj_i1(Co13_C121),
             .Ck_j0(Co14_C130), .Ck_j1(Co14_C131), .Cm_i(C15_C110),
             .Cm_k0(Co15_C140), .Cm_k1(Co15_C141) );
cary_gen I106 ( .C_i(Co8_C71), .Cj_i0(Co9_C80), .Cj_i1(Co9_C81),
             .Ck_j0(Co10_C90), .Ck_j1(Co10_C91), .Cm_i(C11_C71),
             .Cm_k0(Co11_C100), .Cm_k1(Co11_C101) );
cary_gen I107 ( .C_i(Co8_C70), .Cj_i0(Co9_C80), .Cj_i1(Co9_C81),
             .Ck_j0(Co10_C90), .Ck_j1(Co10_C91), .Cm_i(C11_C70),
             .Cm_k0(Co11_C100), .Cm_k1(Co11_C101) );
cary_gen I108 ( .C_i(C19_C151), .Cj_i0(C23_C190), .Cj_i1(C23_C191),
             .Ck_j0(C27_C230), .Ck_j1(C27_C231), .Cm_i(C31_C161),
             .Cm_k0(C31_C270), .Cm_k1(C31_C271) );
cary_gen I109 ( .C_i(C19_C150), .Cj_i0(C23_C190), .Cj_i1(C23_C191),
             .Ck_j0(C27_C230), .Ck_j1(C27_C231), .Cm_i(C31_C160),
             .Cm_k0(C31_C270), .Cm_k1(C31_C271) );
cary_gen I110 ( .C_i(Co28_C271), .Cj_i0(Co29_C280), .Cj_i1(Co29_C281),
             .Ck_j0(Co30_C290), .Ck_j1(Co30_C291), .Cm_i(C31_C271),
             .Cm_k0(Co31_C300), .Cm_k1(Co31_C301) );
cary_gen I111 ( .C_i(Co28_C270), .Cj_i0(Co29_C280), .Cj_i1(Co29_C281),
             .Ck_j0(Co30_C290), .Ck_j1(Co30_C291), .Cm_i(C31_C270),
             .Cm_k0(Co31_C300), .Cm_k1(Co31_C301) );
cary_gen I112 ( .C_i(Co24_C231), .Cj_i0(Co25_C240), .Cj_i1(Co25_C241),
             .Ck_j0(Co26_C250), .Ck_j1(Co26_C251), .Cm_i(C27_C231),
             .Cm_k0(Co27_C260), .Cm_k1(Co27_C261) );
cary_gen I113 ( .C_i(Co24_C230), .Cj_i0(Co25_C240), .Cj_i1(Co25_C241),
             .Ck_j0(Co26_C250), .Ck_j1(Co26_C251), .Cm_i(C27_C230),
             .Cm_k0(Co27_C260), .Cm_k1(Co27_C261) );
cary_gen I114 ( .C_i(Carry3), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
             .Ck_j1(C11_C71), .Cm_i(Carry15b), .Cm_k0(C15_C110),
             .Cm_k1(C15_C111) );
cary_gen I115 ( .C_i(Carry3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
             .Ck_j1(C11_C71), .Cm_i(Carry15a), .Cm_k0(C15_C110),
             .Cm_k1(C15_C111) );
cary_gen I116 ( .C_i(Carry3), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
             .Ck_j1(C11_C71), .Cm_i(Carry15), .Cm_k0(C15_C110),
             .Cm_k1(C15_C111) );
cary_gen I117 ( .C_i(Co20_C191), .Cj_i0(Co21_C200), .Cj_i1(Co21_C201),
             .Ck_j0(Co22_C210), .Ck_j1(Co22_C211), .Cm_i(C23_C191),
             .Cm_k0(Co23_C220), .Cm_k1(Co23_C221) );
cary_gen I118 ( .C_i(Co20_C190), .Cj_i0(Co21_C200), .Cj_i1(Co21_C201),
             .Ck_j0(Co22_C210), .Ck_j1(Co22_C211), .Cm_i(C23_C190),
             .Cm_k0(Co23_C220), .Cm_k1(Co23_C221) );
cary_gen I119 ( .C_i(Co16_C151), .Cj_i0(Co17_C160), .Cj_i1(Co17_C161),
             .Ck_j0(Co18_C170), .Ck_j1(Co18_C171), .Cm_i(C19_C151),
             .Cm_k0(Co19_C180), .Cm_k1(Co19_C181) );
cary_gen I120 ( .C_i(Co16_C150), .Cj_i0(Co17_C160), .Cj_i1(Co17_C161),
             .Ck_j0(Co18_C170), .Ck_j1(Co18_C171), .Cm_i(C19_C150),
             .Cm_k0(Co19_C180), .Cm_k1(Co19_C181) );
cary_gen I121 ( .C_i(Co4_C31), .Cj_i0(Co5_C40), .Cj_i1(Co5_C41), .Ck_j0(Co6_C50),
             .Ck_j1(Co6_C51), .Cm_i(C7_C31), .Cm_k0(Co7_C60), .Cm_k1(Co7_C61) );
cary_gen I122 ( .C_i(Co4_C30), .Cj_i0(Co5_C40), .Cj_i1(Co5_C41), .Ck_j0(Co6_C50),
             .Ck_j1(Co6_C51), .Cm_i(C7_C30), .Cm_k0(Co7_C60), .Cm_k1(Co7_C61) );

endmodule // borrow32

`endif

`ifdef borrow16
`else
`define borrow16
module borrow16( a , b, Borrow3, Bo, C11_C70, C11_C71, C7_C30, C7_C31, Co0_Ci0,
                 Co0_Ci1, Co10_C90, Co10_C91, Co12_C110, Co12_C111, Co13_C120,
                 Co13_C121, Co14_C130, Co14_C131, Co1_C00, Co1_C01, Co2_C10,
                 Co2_C11, Co3_C20, Co3_C21, Co4_C30, Co4_C31, Co5_C40,
                 Co5_C41, Co6_C50, Co6_C51, Co8_C70, Co8_C71, Co9_C80,
                 Co9_C81, D );
 input [15:0] a;
 input [15:0] b;
output Bo;
input Borrow3;
output C11_C70, C11_C71, C7_C30, C7_C31, Co0_Ci0, Co0_Ci1, Co10_C90, Co10_C91,
Co12_C110, Co12_C111, Co13_C120, Co13_C121, Co14_C130, Co14_C131,
Co1_C00, Co1_C01, Co2_C10, Co2_C11, Co3_C20, Co3_C21, Co4_C30, Co4_C31,
Co5_C40, Co5_C41, Co6_C50, Co6_C51, Co8_C70, Co8_C71, Co9_C80, Co9_C81;
 output [15:0] D;
wire Co7_C60;
wire Co7_C61;
wire Co11_C100;
wire Co11_C101;
wire Co15_C140;
wire Co15_C141;
wire C15_C110;
wire C15_C111;

dif_b0 I_107 ( .Ax(a[0]), .Bo_Bi0(Co0_Ci0), .Bo_Bi1(Co0_Ci1), .Bx(b[0]) );
bo_gen I111 ( .C_i(Borrow3), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
           .Ck_j1(C11_C71), .Cm_i(Bo), .Cm_k0(C15_C110), .Cm_k1(C15_C111) );
dif_b I_105 ( .Ax(a[1]), .Bo_Bi0(Co1_C00), .Bo_Bi1(Co1_C01), .Bx(b[1]),
           .Sub_Dif(D[1]) );
dif_b I_103 ( .Ax(a[2]), .Bo_Bi0(Co2_C10), .Bo_Bi1(Co2_C11), .Bx(b[2]),
           .Sub_Dif(D[2]) );
dif_b I_102 ( .Ax(a[3]), .Bo_Bi0(Co3_C20), .Bo_Bi1(Co3_C21), .Bx(b[3]),
           .Sub_Dif(D[3]) );
dif_b I_101 ( .Ax(a[4]), .Bo_Bi0(Co4_C30), .Bo_Bi1(Co4_C31), .Bx(b[4]),
           .Sub_Dif(D[4]) );
dif_b I_100 ( .Ax(a[5]), .Bo_Bi0(Co5_C40), .Bo_Bi1(Co5_C41), .Bx(b[5]),
           .Sub_Dif(D[5]) );
dif_b I_99 ( .Ax(a[6]), .Bo_Bi0(Co6_C50), .Bo_Bi1(Co6_C51), .Bx(b[6]),
          .Sub_Dif(D[6]) );
dif_b I_98 ( .Ax(a[7]), .Bo_Bi0(Co7_C60), .Bo_Bi1(Co7_C61), .Bx(b[7]),
          .Sub_Dif(D[7]) );
dif_b I_97 ( .Ax(a[8]), .Bo_Bi0(Co8_C70), .Bo_Bi1(Co8_C71), .Bx(b[8]),
          .Sub_Dif(D[8]) );
dif_b I_96 ( .Ax(a[9]), .Bo_Bi0(Co9_C80), .Bo_Bi1(Co9_C81), .Bx(b[9]),
          .Sub_Dif(D[9]) );
dif_b I_95 ( .Ax(a[10]), .Bo_Bi0(Co10_C90), .Bo_Bi1(Co10_C91), .Bx(b[10]),
          .Sub_Dif(D[10]) );
dif_b I_94 ( .Ax(a[11]), .Bo_Bi0(Co11_C100), .Bo_Bi1(Co11_C101), .Bx(b[11]),
          .Sub_Dif(D[11]) );
dif_b I_93 ( .Ax(a[12]), .Bo_Bi0(Co12_C110), .Bo_Bi1(Co12_C111), .Bx(b[12]),
          .Sub_Dif(D[12]) );
dif_b I_91 ( .Ax(a[14]), .Bo_Bi0(Co14_C130), .Bo_Bi1(Co14_C131), .Bx(b[14]),
          .Sub_Dif(D[14]) );
dif_b I_90 ( .Ax(a[15]), .Bo_Bi0(Co15_C140), .Bo_Bi1(Co15_C141), .Bx(b[15]),
          .Sub_Dif(D[15]) );
dif_b I_92 ( .Ax(a[13]), .Bo_Bi0(Co13_C120), .Bo_Bi1(Co13_C121), .Bx(b[13]),
          .Sub_Dif(D[13]) );
cary_gen I105 ( .C_i(Co12_C111), .Cj_i0(Co13_C120), .Cj_i1(Co13_C121),
             .Ck_j0(Co14_C130), .Ck_j1(Co14_C131), .Cm_i(C15_C111),
             .Cm_k0(Co15_C140), .Cm_k1(Co15_C141) );
cary_gen I106 ( .C_i(Co12_C110), .Cj_i0(Co13_C120), .Cj_i1(Co13_C121),
             .Ck_j0(Co14_C130), .Ck_j1(Co14_C131), .Cm_i(C15_C110),
             .Cm_k0(Co15_C140), .Cm_k1(Co15_C141) );
cary_gen I107 ( .C_i(Co8_C71), .Cj_i0(Co9_C80), .Cj_i1(Co9_C81),
             .Ck_j0(Co10_C90), .Ck_j1(Co10_C91), .Cm_i(C11_C71),
             .Cm_k0(Co11_C100), .Cm_k1(Co11_C101) );
cary_gen I108 ( .C_i(Co8_C70), .Cj_i0(Co9_C80), .Cj_i1(Co9_C81),
             .Ck_j0(Co10_C90), .Ck_j1(Co10_C91), .Cm_i(C11_C70),
             .Cm_k0(Co11_C100), .Cm_k1(Co11_C101) );
cary_gen I109 ( .C_i(Co4_C31), .Cj_i0(Co5_C40), .Cj_i1(Co5_C41), .Ck_j0(Co6_C50),
             .Ck_j1(Co6_C51), .Cm_i(C7_C31), .Cm_k0(Co7_C60), .Cm_k1(Co7_C61) );
cary_gen I110 ( .C_i(Co4_C30), .Cj_i0(Co5_C40), .Cj_i1(Co5_C41), .Ck_j0(Co6_C50),
             .Ck_j1(Co6_C51), .Cm_i(C7_C30), .Cm_k0(Co7_C60), .Cm_k1(Co7_C61) );

endmodule // borrow16

`endif

`ifdef dif16
`else
`define dif16
module dif16( a , b, Bin, C11_C70, C11_C71, C7_C30, C7_C31, Co0_Ci0, Co0_Ci1,
              Co10_C90, Co10_C91, Co12_C110, Co12_C111, Co13_C120, Co13_C121,
              Co14_C130, Co14_C131, Co1_C00, Co1_C01, Co2_C10, Co2_C11,
              Co3_C20, Co3_C21, Co4_C30, Co4_C31, Co5_C40, Co5_C41, Co6_C50,
              Co6_C51, Co8_C70, Co8_C71, Co9_C80, Co9_C81, D, Borrow3, Diffi );
 input [0:0] a;
 input [0:0] b;
input Bin;
output Borrow3;
input C11_C70, C11_C71, C7_C30, C7_C31, Co0_Ci0, Co0_Ci1, Co10_C90, Co10_C91,
Co12_C110, Co12_C111, Co13_C120, Co13_C121, Co14_C130, Co14_C131,
Co1_C00, Co1_C01, Co2_C10, Co2_C11, Co3_C20, Co3_C21, Co4_C30, Co4_C31,
Co5_C40, Co5_C41, Co6_C50, Co6_C51, Co8_C70, Co8_C71, Co9_C80, Co9_C81;
 input [15:0] D;
 output [15:0] Diffi;
wire Borrow_0;
wire Borrow3a;
wire N_189;
wire N_190;
wire N_191;
wire N_192;
wire N_193;
wire N_194;
wire N_195;
wire N_196;
wire N_197;
wire N_198;
wire N_199;
wire N_200;
supply0 gnd;

borrow0 I_135 ( .A(a[0]), .B(b[0]), .Bin(Bin), .Bout(Borrow_0) );
dif0 I_134 ( .A(a[0]), .B(b[0]), .Bin(Bin), .d0(Diffi[0]) );
sum2_gen I150 ( .C_i(Borrow3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
             .Ck_j1(C11_C71), .Sk_0(N_200), .Sk_1(N_197), .Sk_i(Diffi[15]) );
sum2_gen I151 ( .C_i(Borrow3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
             .Ck_j1(C11_C71), .Sk_0(N_198), .Sk_1(N_196), .Sk_i(Diffi[14]) );
sum2_gen I152 ( .C_i(Borrow3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
             .Ck_j1(C11_C71), .Sk_0(N_199), .Sk_1(N_195), .Sk_i(Diffi[13]) );
sum2_gen I140 ( .C_i(gnd), .Cj_i0(Borrow3a), .Cj_i1(gnd), .Ck_j0(C7_C30),
             .Ck_j1(C7_C31), .Sk_0(N_194), .Sk_1(N_191), .Sk_i(Diffi[11]) );
sum2_gen I141 ( .C_i(gnd), .Cj_i0(Borrow3a), .Cj_i1(gnd), .Ck_j0(C7_C30),
             .Ck_j1(C7_C31), .Sk_0(N_192), .Sk_1(N_193), .Sk_i(Diffi[10]) );
sum2_gen I134 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Borrow3), .Ck_j1(gnd),
             .Sk_0(N_189), .Sk_1(N_190), .Sk_i(Diffi[7]) );
cary_gen I148 ( .C_i(Borrow_0), .Cj_i0(Co1_C00), .Cj_i1(Co1_C01),
             .Ck_j0(Co2_C10), .Ck_j1(Co2_C11), .Cm_i(Borrow3a),
             .Cm_k0(Co3_C20), .Cm_k1(Co3_C21) );
cary_gen I149 ( .C_i(Borrow_0), .Cj_i0(Co1_C00), .Cj_i1(Co1_C01),
             .Ck_j0(Co2_C10), .Ck_j1(Co2_C11), .Cm_i(Borrow3),
             .Cm_k0(Co3_C20), .Cm_k1(Co3_C21) );
sum_gen I153 ( .C_i(Co12_C111), .Cj_i0(Co13_C120), .Cj_i1(Co13_C121),
            .Ck_j0(Co14_C130), .Ck_j1(Co14_C131), .Sk_01(D[15]), .Sk_i(N_197) );
sum_gen I154 ( .C_i(Co12_C110), .Cj_i0(Co13_C120), .Cj_i1(Co13_C121),
            .Ck_j0(Co14_C130), .Ck_j1(Co14_C131), .Sk_01(D[15]), .Sk_i(N_200) );
sum_gen I155 ( .C_i(gnd), .Cj_i0(Co12_C111), .Cj_i1(gnd), .Ck_j0(Co13_C120),
            .Ck_j1(Co13_C121), .Sk_01(D[14]), .Sk_i(N_196) );
sum_gen I156 ( .C_i(gnd), .Cj_i0(Co12_C110), .Cj_i1(gnd), .Ck_j0(Co13_C120),
            .Ck_j1(Co13_C121), .Sk_01(D[14]), .Sk_i(N_198) );
sum_gen I157 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Co12_C111),
            .Ck_j1(gnd), .Sk_01(D[13]), .Sk_i(N_195) );
sum_gen I158 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Co12_C110),
            .Ck_j1(gnd), .Sk_01(D[13]), .Sk_i(N_199) );
sum_gen I159 ( .C_i(Borrow3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
            .Ck_j1(C11_C71), .Sk_01(D[12]), .Sk_i(Diffi[12]) );
sum_gen I142 ( .C_i(Co8_C71), .Cj_i0(Co9_C80), .Cj_i1(Co9_C81), .Ck_j0(Co10_C90),
            .Ck_j1(Co10_C91), .Sk_01(D[11]), .Sk_i(N_191) );
sum_gen I143 ( .C_i(Co8_C70), .Cj_i0(Co9_C80), .Cj_i1(Co9_C81), .Ck_j0(Co10_C90),
            .Ck_j1(Co10_C91), .Sk_01(D[11]), .Sk_i(N_194) );
sum_gen I144 ( .C_i(gnd), .Cj_i0(Co8_C71), .Cj_i1(gnd), .Ck_j0(Co9_C80),
            .Ck_j1(Co9_C81), .Sk_01(D[10]), .Sk_i(N_193) );
sum_gen I145 ( .C_i(gnd), .Cj_i0(Co8_C70), .Cj_i1(gnd), .Ck_j0(Co9_C80),
            .Ck_j1(Co9_C81), .Sk_01(D[10]), .Sk_i(N_192) );
sum_gen I146 ( .C_i(Borrow3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(Co8_C70),
            .Ck_j1(Co8_C71), .Sk_01(D[9]), .Sk_i(Diffi[9]) );
sum_gen I147 ( .C_i(gnd), .Cj_i0(Borrow3a), .Cj_i1(gnd), .Ck_j0(C7_C30),
            .Ck_j1(C7_C31), .Sk_01(D[8]), .Sk_i(Diffi[8]) );
sum_gen I135 ( .C_i(Co4_C31), .Cj_i0(Co5_C40), .Cj_i1(Co5_C41), .Ck_j0(Co6_C50),
            .Ck_j1(Co6_C51), .Sk_01(D[7]), .Sk_i(N_190) );
sum_gen I136 ( .C_i(Co4_C30), .Cj_i0(Co5_C40), .Cj_i1(Co5_C41), .Ck_j0(Co6_C50),
            .Ck_j1(Co6_C51), .Sk_01(D[7]), .Sk_i(N_189) );
sum_gen I137 ( .C_i(Borrow3), .Cj_i0(Co4_C30), .Cj_i1(Co4_C31), .Ck_j0(Co5_C40),
            .Ck_j1(Co5_C41), .Sk_01(D[6]), .Sk_i(Diffi[6]) );
sum_gen I138 ( .C_i(gnd), .Cj_i0(Borrow3), .Cj_i1(gnd), .Ck_j0(Co4_C30),
            .Ck_j1(Co4_C31), .Sk_01(D[5]), .Sk_i(Diffi[5]) );
sum_gen I139 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Borrow3), .Ck_j1(gnd),
            .Sk_01(D[4]), .Sk_i(Diffi[4]) );
sum_gen I131 ( .C_i(Borrow_0), .Cj_i0(Co1_C00), .Cj_i1(Co1_C01), .Ck_j0(Co2_C10),
            .Ck_j1(Co2_C11), .Sk_01(D[3]), .Sk_i(Diffi[3]) );
sum_gen I132 ( .C_i(Bin), .Cj_i0(Co0_Ci1), .Cj_i1(Co0_Ci0), .Ck_j0(Co1_C00),
            .Ck_j1(Co1_C01), .Sk_01(D[2]), .Sk_i(Diffi[2]) );
sum_gen I133 ( .C_i(gnd), .Cj_i0(Bin), .Cj_i1(gnd), .Ck_j0(Co0_Ci1),
            .Ck_j1(Co0_Ci0), .Sk_01(D[1]), .Sk_i(Diffi[1]) );

endmodule // dif16

`endif

`ifdef carry32
`else
`define carry32
module carry32( a , b, Carry3, Carry3a, C11_C70, C11_C71, C19_C150, C19_C151,
                C23_C190, C23_C191, C27_C230, C27_C231, C7_C30, C7_C31,
                Carry15, Carry15a, Carry15b, Co, Co0_Ci0, Co0_Ci1, Co10_C90,
                Co10_C91, Co12_C110, Co12_C111, Co13_C120, Co13_C121,
                Co14_C130, Co14_C131, Co16_C150, Co16_C151, Co17_C160,
                Co17_C161, Co18_C170, Co18_C171, Co1_C00, Co1_C01, Co20_C190,
                Co20_C191, Co21_C200, Co21_C201, Co22_C210, Co22_C211,
                Co24_C230, Co24_C231, Co25_C240, Co25_C241, Co26_C250,
                Co26_C251, Co28_C270, Co28_C271, Co29_C280, Co29_C281,
                Co2_C10, Co2_C11, Co30_C290, Co30_C291, Co3_C20, Co3_C21,
                Co4_C30, Co4_C31, Co5_C40, Co5_C41, Co6_C50, Co6_C51, Co8_C70,
                Co8_C71, Co9_C80, Co9_C81, S );
 input [31:0] a;
 input [31:0] b;
output C11_C70, C11_C71, C19_C150, C19_C151, C23_C190, C23_C191, C27_C230,
C27_C231, C7_C30, C7_C31, Carry15, Carry15a, Carry15b;
input Carry3, Carry3a;
output Co, Co0_Ci0, Co0_Ci1, Co10_C90, Co10_C91, Co12_C110, Co12_C111,
Co13_C120, Co13_C121, Co14_C130, Co14_C131, Co16_C150, Co16_C151,
Co17_C160, Co17_C161, Co18_C170, Co18_C171, Co1_C00, Co1_C01,
Co20_C190, Co20_C191, Co21_C200, Co21_C201, Co22_C210, Co22_C211,
Co24_C230, Co24_C231, Co25_C240, Co25_C241, Co26_C250, Co26_C251,
Co28_C270, Co28_C271, Co29_C280, Co29_C281, Co2_C10, Co2_C11,
Co30_C290, Co30_C291, Co3_C20, Co3_C21, Co4_C30, Co4_C31, Co5_C40,
Co5_C41, Co6_C50, Co6_C51, Co8_C70, Co8_C71, Co9_C80, Co9_C81;
 output [31:0] S;
supply0 gnd;
wire C31_C160;
wire C31_C161;
wire Co19_C180;
wire Co19_C181;
wire Co23_C220;
wire Co23_C221;
wire Co7_C60;
wire Co7_C61;
wire Co11_C100;
wire Co11_C101;
wire Co15_C140;
wire Co15_C141;
wire Co27_C260;
wire Co27_C261;
wire Co31_C300;
wire Co31_C301;
wire C31_C270;
wire C31_C271;
wire C15_C110;
wire C15_C111;

sum_c0 I_74 ( .Ax(a[0]), .Bx(b[0]), .Co_Ci0(Co0_Ci0), .Co_Ci1(Co0_Ci1) );
cary_gen I86 ( .C_i(Carry3), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
            .Ck_j1(C11_C71), .Cm_i(Carry15), .Cm_k0(C15_C110),
            .Cm_k1(C15_C111) );
cary_gen I87 ( .C_i(Carry3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
            .Ck_j1(C11_C71), .Cm_i(Carry15a), .Cm_k0(C15_C110),
            .Cm_k1(C15_C111) );
cary_gen I88 ( .C_i(Carry3), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
            .Ck_j1(C11_C71), .Cm_i(Carry15b), .Cm_k0(C15_C110),
            .Cm_k1(C15_C111) );
cary_gen I89 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Carry15), .Ck_j1(gnd),
            .Cm_i(Co), .Cm_k0(C31_C160), .Cm_k1(C31_C161) );
cary_gen I90 ( .C_i(C19_C151), .Cj_i0(C23_C190), .Cj_i1(C23_C191),
            .Ck_j0(C27_C230), .Ck_j1(C27_C231), .Cm_i(C31_C161),
            .Cm_k0(C31_C270), .Cm_k1(C31_C271) );
cary_gen I91 ( .C_i(C19_C150), .Cj_i0(C23_C190), .Cj_i1(C23_C191),
            .Ck_j0(C27_C230), .Ck_j1(C27_C231), .Cm_i(C31_C160),
            .Cm_k0(C31_C270), .Cm_k1(C31_C271) );
cary_gen I82 ( .C_i(Co28_C271), .Cj_i0(Co29_C280), .Cj_i1(Co29_C281),
            .Ck_j0(Co30_C290), .Ck_j1(Co30_C291), .Cm_i(C31_C271),
            .Cm_k0(Co31_C300), .Cm_k1(Co31_C301) );
cary_gen I83 ( .C_i(Co28_C270), .Cj_i0(Co29_C280), .Cj_i1(Co29_C281),
            .Ck_j0(Co30_C290), .Ck_j1(Co30_C291), .Cm_i(C31_C270),
            .Cm_k0(Co31_C300), .Cm_k1(Co31_C301) );
cary_gen I84 ( .C_i(Co24_C231), .Cj_i0(Co25_C240), .Cj_i1(Co25_C241),
            .Ck_j0(Co26_C250), .Ck_j1(Co26_C251), .Cm_i(C27_C231),
            .Cm_k0(Co27_C260), .Cm_k1(Co27_C261) );
cary_gen I85 ( .C_i(Co24_C230), .Cj_i0(Co25_C240), .Cj_i1(Co25_C241),
            .Ck_j0(Co26_C250), .Ck_j1(Co26_C251), .Cm_i(C27_C230),
            .Cm_k0(Co27_C260), .Cm_k1(Co27_C261) );
cary_gen I76 ( .C_i(Co20_C191), .Cj_i0(Co21_C200), .Cj_i1(Co21_C201),
            .Ck_j0(Co22_C210), .Ck_j1(Co22_C211), .Cm_i(C23_C191),
            .Cm_k0(Co23_C220), .Cm_k1(Co23_C221) );
cary_gen I77 ( .C_i(Co20_C190), .Cj_i0(Co21_C200), .Cj_i1(Co21_C201),
            .Ck_j0(Co22_C210), .Ck_j1(Co22_C211), .Cm_i(C23_C190),
            .Cm_k0(Co23_C220), .Cm_k1(Co23_C221) );
cary_gen I78 ( .C_i(Co16_C151), .Cj_i0(Co17_C160), .Cj_i1(Co17_C161),
            .Ck_j0(Co18_C170), .Ck_j1(Co18_C171), .Cm_i(C19_C151),
            .Cm_k0(Co19_C180), .Cm_k1(Co19_C181) );
cary_gen I79 ( .C_i(Co16_C150), .Cj_i0(Co17_C160), .Cj_i1(Co17_C161),
            .Ck_j0(Co18_C170), .Ck_j1(Co18_C171), .Cm_i(C19_C150),
            .Cm_k0(Co19_C180), .Cm_k1(Co19_C181) );
cary_gen I80 ( .C_i(Co12_C111), .Cj_i0(Co13_C120), .Cj_i1(Co13_C121),
            .Ck_j0(Co14_C130), .Ck_j1(Co14_C131), .Cm_i(C15_C111),
            .Cm_k0(Co15_C140), .Cm_k1(Co15_C141) );
cary_gen I81 ( .C_i(Co12_C110), .Cj_i0(Co13_C120), .Cj_i1(Co13_C121),
            .Ck_j0(Co14_C130), .Ck_j1(Co14_C131), .Cm_i(C15_C110),
            .Cm_k0(Co15_C140), .Cm_k1(Co15_C141) );
cary_gen I72 ( .C_i(Co8_C71), .Cj_i0(Co9_C80), .Cj_i1(Co9_C81), .Ck_j0(Co10_C90),
            .Ck_j1(Co10_C91), .Cm_i(C11_C71), .Cm_k0(Co11_C100),
            .Cm_k1(Co11_C101) );
cary_gen I73 ( .C_i(Co8_C70), .Cj_i0(Co9_C80), .Cj_i1(Co9_C81), .Ck_j0(Co10_C90),
            .Ck_j1(Co10_C91), .Cm_i(C11_C70), .Cm_k0(Co11_C100),
            .Cm_k1(Co11_C101) );
cary_gen I74 ( .C_i(Co4_C31), .Cj_i0(Co5_C40), .Cj_i1(Co5_C41), .Ck_j0(Co6_C50),
            .Ck_j1(Co6_C51), .Cm_i(C7_C31), .Cm_k0(Co7_C60), .Cm_k1(Co7_C61) );
cary_gen I75 ( .C_i(Co4_C30), .Cj_i0(Co5_C40), .Cj_i1(Co5_C41), .Ck_j0(Co6_C50),
            .Ck_j1(Co6_C51), .Cm_i(C7_C30), .Cm_k0(Co7_C60), .Cm_k1(Co7_C61) );
sum_c I_45 ( .Ax(a[16]), .Bx(b[16]), .Co_Ci0(Co16_C150), .Co_Ci1(Co16_C151),
          .Sub_Sum(S[16]) );
sum_c I_46 ( .Ax(a[17]), .Bx(b[17]), .Co_Ci0(Co17_C160), .Co_Ci1(Co17_C161),
          .Sub_Sum(S[17]) );
sum_c I_48 ( .Ax(a[19]), .Bx(b[19]), .Co_Ci0(Co19_C180), .Co_Ci1(Co19_C181),
          .Sub_Sum(S[19]) );
sum_c I_47 ( .Ax(a[18]), .Bx(b[18]), .Co_Ci0(Co18_C170), .Co_Ci1(Co18_C171),
          .Sub_Sum(S[18]) );
sum_c I_49 ( .Ax(a[20]), .Bx(b[20]), .Co_Ci0(Co20_C190), .Co_Ci1(Co20_C191),
          .Sub_Sum(S[20]) );
sum_c I_50 ( .Ax(a[21]), .Bx(b[21]), .Co_Ci0(Co21_C200), .Co_Ci1(Co21_C201),
          .Sub_Sum(S[21]) );
sum_c I_51 ( .Ax(a[22]), .Bx(b[22]), .Co_Ci0(Co22_C210), .Co_Ci1(Co22_C211),
          .Sub_Sum(S[22]) );
sum_c I_52 ( .Ax(a[23]), .Bx(b[23]), .Co_Ci0(Co23_C220), .Co_Ci1(Co23_C221),
          .Sub_Sum(S[23]) );
sum_c I_53 ( .Ax(a[24]), .Bx(b[24]), .Co_Ci0(Co24_C230), .Co_Ci1(Co24_C231),
          .Sub_Sum(S[24]) );
sum_c I_54 ( .Ax(a[25]), .Bx(b[25]), .Co_Ci0(Co25_C240), .Co_Ci1(Co25_C241),
          .Sub_Sum(S[25]) );
sum_c I_55 ( .Ax(a[26]), .Bx(b[26]), .Co_Ci0(Co26_C250), .Co_Ci1(Co26_C251),
          .Sub_Sum(S[26]) );
sum_c I_56 ( .Ax(a[27]), .Bx(b[27]), .Co_Ci0(Co27_C260), .Co_Ci1(Co27_C261),
          .Sub_Sum(S[27]) );
sum_c I_57 ( .Ax(a[28]), .Bx(b[28]), .Co_Ci0(Co28_C270), .Co_Ci1(Co28_C271),
          .Sub_Sum(S[28]) );
sum_c I_58 ( .Ax(a[29]), .Bx(b[29]), .Co_Ci0(Co29_C280), .Co_Ci1(Co29_C281),
          .Sub_Sum(S[29]) );
sum_c I_59 ( .Ax(a[30]), .Bx(b[30]), .Co_Ci0(Co30_C290), .Co_Ci1(Co30_C291),
          .Sub_Sum(S[30]) );
sum_c I_44 ( .Ax(a[31]), .Bx(b[31]), .Co_Ci0(Co31_C300), .Co_Ci1(Co31_C301),
          .Sub_Sum(S[31]) );
sum_c s1 ( .Ax(a[1]), .Bx(b[1]), .Co_Ci0(Co1_C00), .Co_Ci1(Co1_C01),
        .Sub_Sum(S[1]) );
sum_c s2 ( .Ax(a[2]), .Bx(b[2]), .Co_Ci0(Co2_C10), .Co_Ci1(Co2_C11),
        .Sub_Sum(S[2]) );
sum_c s3 ( .Ax(a[3]), .Bx(b[3]), .Co_Ci0(Co3_C20), .Co_Ci1(Co3_C21),
        .Sub_Sum(S[3]) );
sum_c s4 ( .Ax(a[4]), .Bx(b[4]), .Co_Ci0(Co4_C30), .Co_Ci1(Co4_C31),
        .Sub_Sum(S[4]) );
sum_c s5 ( .Ax(a[5]), .Bx(b[5]), .Co_Ci0(Co5_C40), .Co_Ci1(Co5_C41),
        .Sub_Sum(S[5]) );
sum_c s6 ( .Ax(a[6]), .Bx(b[6]), .Co_Ci0(Co6_C50), .Co_Ci1(Co6_C51),
        .Sub_Sum(S[6]) );
sum_c s7 ( .Ax(a[7]), .Bx(b[7]), .Co_Ci0(Co7_C60), .Co_Ci1(Co7_C61),
        .Sub_Sum(S[7]) );
sum_c s8 ( .Ax(a[8]), .Bx(b[8]), .Co_Ci0(Co8_C70), .Co_Ci1(Co8_C71),
        .Sub_Sum(S[8]) );
sum_c s9 ( .Ax(a[9]), .Bx(b[9]), .Co_Ci0(Co9_C80), .Co_Ci1(Co9_C81),
        .Sub_Sum(S[9]) );
sum_c s10 ( .Ax(a[10]), .Bx(b[10]), .Co_Ci0(Co10_C90), .Co_Ci1(Co10_C91),
         .Sub_Sum(S[10]) );
sum_c s11 ( .Ax(a[11]), .Bx(b[11]), .Co_Ci0(Co11_C100), .Co_Ci1(Co11_C101),
         .Sub_Sum(S[11]) );
sum_c s12 ( .Ax(a[12]), .Bx(b[12]), .Co_Ci0(Co12_C110), .Co_Ci1(Co12_C111),
         .Sub_Sum(S[12]) );
sum_c s13 ( .Ax(a[13]), .Bx(b[13]), .Co_Ci0(Co13_C120), .Co_Ci1(Co13_C121),
         .Sub_Sum(S[13]) );
sum_c s14 ( .Ax(a[14]), .Bx(b[14]), .Co_Ci0(Co14_C130), .Co_Ci1(Co14_C131),
         .Sub_Sum(S[14]) );
sum_c s15 ( .Ax(a[15]), .Bx(b[15]), .Co_Ci0(Co15_C140), .Co_Ci1(Co15_C141),
         .Sub_Sum(S[15]) );

endmodule // carry32

`endif

`ifdef sum32
`else
`define sum32
module sum32( a , b, C11_C70, C11_C71, C19_C150, C19_C151, C23_C190, C23_C191,
              C27_C230, C27_C231, C7_C30, C7_C31, Carry15, Carry15a, Carry15b,
              Cin, Co0_Ci0, Co0_Ci1, Co10_C90, Co10_C91, Co12_C110, Co12_C111,
              Co13_C120, Co13_C121, Co14_C130, Co14_C131, Co16_C150,
              Co16_C151, Co17_C160, Co17_C161, Co18_C170, Co18_C171, Co1_C00,
              Co1_C01, Co20_C190, Co20_C191, Co21_C200, Co21_C201, Co22_C210,
              Co22_C211, Co24_C230, Co24_C231, Co25_C240, Co25_C241,
              Co26_C250, Co26_C251, Co28_C270, Co28_C271, Co29_C280,
              Co29_C281, Co2_C10, Co2_C11, Co30_C290, Co30_C291, Co3_C20,
              Co3_C21, Co4_C30, Co4_C31, Co5_C40, Co5_C41, Co6_C50, Co6_C51,
              Co8_C70, Co8_C71, Co9_C80, Co9_C81, S, Carry3, Carry3a, Sumi );
 input [0:0] a;
 input [0:0] b;
input C11_C70, C11_C71, C19_C150, C19_C151, C23_C190, C23_C191, C27_C230,
C27_C231, C7_C30, C7_C31, Carry15, Carry15a, Carry15b;
output Carry3, Carry3a;
input Cin, Co0_Ci0, Co0_Ci1, Co10_C90, Co10_C91, Co12_C110, Co12_C111,
Co13_C120, Co13_C121, Co14_C130, Co14_C131, Co16_C150, Co16_C151,
Co17_C160, Co17_C161, Co18_C170, Co18_C171, Co1_C00, Co1_C01,
Co20_C190, Co20_C191, Co21_C200, Co21_C201, Co22_C210, Co22_C211,
Co24_C230, Co24_C231, Co25_C240, Co25_C241, Co26_C250, Co26_C251,
Co28_C270, Co28_C271, Co29_C280, Co29_C281, Co2_C10, Co2_C11,
Co30_C290, Co30_C291, Co3_C20, Co3_C21, Co4_C30, Co4_C31, Co5_C40,
Co5_C41, Co6_C50, Co6_C51, Co8_C70, Co8_C71, Co9_C80, Co9_C81;
 input [31:0] S;
 output [31:0] Sumi;
wire Carry_0;
wire N_233;
wire N_234;
wire N_227;
wire N_228;
wire N_229;
wire N_230;
wire N_231;
wire N_232;
wire N_213;
wire N_214;
wire N_215;
wire N_216;
wire N_217;
wire N_218;
wire N_219;
wire N_220;
wire N_221;
wire N_222;
wire N_223;
wire N_224;
wire N_225;
wire N_226;
wire N_207;
wire N_208;
wire N_209;
wire N_210;
wire N_211;
wire N_212;
wire N_201;
wire N_202;
wire N_203;
wire N_204;
wire N_205;
wire N_206;
supply0 gnd;

mux2x0 I_133 ( .A(N_221), .B(N_222), .Q(Sumi[31]), .S(Carry15b) );
sum2_gen I162 ( .C_i(gnd), .Cj_i0(Carry15), .Cj_i1(gnd), .Ck_j0(C19_C150),
             .Ck_j1(C19_C151), .Sk_0(N_226), .Sk_1(N_225), .Sk_i(Sumi[23]) );
sum2_gen I163 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Carry15), .Ck_j1(gnd),
             .Sk_0(N_224), .Sk_1(N_223), .Sk_i(Sumi[22]) );
sum2_gen I164 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Carry15a),
             .Ck_j1(gnd), .Sk_0(N_234), .Sk_1(N_233), .Sk_i(Sumi[19]) );
sum2_gen I165 ( .C_i(Carry15a), .Cj_i0(C19_C150), .Cj_i1(C19_C151),
             .Ck_j0(C23_C190), .Ck_j1(C23_C191), .Sk_0(N_214), .Sk_1(N_213),
             .Sk_i(Sumi[28]) );
sum2_gen I166 ( .C_i(Carry15b), .Cj_i0(C19_C150), .Cj_i1(C19_C151),
             .Ck_j0(C23_C190), .Ck_j1(C23_C191), .Sk_0(N_216), .Sk_1(N_215),
             .Sk_i(Sumi[29]) );
sum2_gen I167 ( .C_i(Carry15b), .Cj_i0(C19_C150), .Cj_i1(C19_C151),
             .Ck_j0(C23_C190), .Ck_j1(C23_C191), .Sk_0(N_218), .Sk_1(N_217),
             .Sk_i(Sumi[30]) );
sum2_gen I168 ( .C_i(C19_C150), .Cj_i0(C23_C190), .Cj_i1(C23_C191),
             .Ck_j0(C27_C230), .Ck_j1(C27_C231), .Sk_0(N_219), .Sk_1(N_220),
             .Sk_i(N_221) );
sum2_gen I169 ( .C_i(C19_C151), .Cj_i0(C23_C190), .Cj_i1(C23_C191),
             .Ck_j0(C27_C230), .Ck_j1(C27_C231), .Sk_0(N_219), .Sk_1(N_220),
             .Sk_i(N_222) );
sum2_gen I170 ( .C_i(Carry15b), .Cj_i0(C19_C150), .Cj_i1(C19_C151),
             .Ck_j0(C23_C190), .Ck_j1(C23_C191), .Sk_0(N_232), .Sk_1(N_231),
             .Sk_i(Sumi[27]) );
sum2_gen I171 ( .C_i(Carry15b), .Cj_i0(C19_C150), .Cj_i1(C19_C151),
             .Ck_j0(C23_C190), .Ck_j1(C23_C191), .Sk_0(N_230), .Sk_1(N_229),
             .Sk_i(Sumi[26]) );
sum2_gen I172 ( .C_i(Carry15b), .Cj_i0(C19_C150), .Cj_i1(C19_C151),
             .Ck_j0(C23_C190), .Ck_j1(C23_C191), .Sk_0(N_228), .Sk_1(N_227),
             .Sk_i(Sumi[25]) );
sum2_gen I159 ( .C_i(Carry3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
             .Ck_j1(C11_C71), .Sk_0(N_212), .Sk_1(N_211), .Sk_i(Sumi[15]) );
sum2_gen I160 ( .C_i(Carry3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
             .Ck_j1(C11_C71), .Sk_0(N_210), .Sk_1(N_209), .Sk_i(Sumi[14]) );
sum2_gen I161 ( .C_i(Carry3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
             .Ck_j1(C11_C71), .Sk_0(N_208), .Sk_1(N_207), .Sk_i(Sumi[13]) );
sum2_gen I156 ( .C_i(gnd), .Cj_i0(Carry3a), .Cj_i1(gnd), .Ck_j0(C7_C30),
             .Ck_j1(C7_C31), .Sk_0(N_202), .Sk_1(N_201), .Sk_i(Sumi[11]) );
sum2_gen I157 ( .C_i(gnd), .Cj_i0(Carry3a), .Cj_i1(gnd), .Ck_j0(C7_C30),
             .Ck_j1(C7_C31), .Sk_0(N_203), .Sk_1(N_204), .Sk_i(Sumi[10]) );
sum2_gen I158 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Carry3), .Ck_j1(gnd),
             .Sk_0(N_205), .Sk_1(N_206), .Sk_i(Sumi[7]) );
cary_gen I133 ( .C_i(Carry_0), .Cj_i0(Co1_C00), .Cj_i1(Co1_C01), .Ck_j0(Co2_C10),
             .Ck_j1(Co2_C11), .Cm_i(Carry3a), .Cm_k0(Co3_C20),
             .Cm_k1(Co3_C21) );
cary_gen I134 ( .C_i(Carry_0), .Cj_i0(Co1_C00), .Cj_i1(Co1_C01), .Ck_j0(Co2_C10),
             .Ck_j1(Co2_C11), .Cm_i(Carry3), .Cm_k0(Co3_C20), .Cm_k1(Co3_C21) );
carry0 I131 ( .A(a[0]), .B(b[0]), .Cin(Cin), .Cout(Carry_0) );
sum_gen I173 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(C27_C230), .Ck_j1(gnd),
            .Sk_01(S[28]), .Sk_i(N_214) );
sum_gen I174 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(C27_C231), .Ck_j1(gnd),
            .Sk_01(S[28]), .Sk_i(N_213) );
sum_gen I175 ( .C_i(Co28_C271), .Cj_i0(Co29_C280), .Cj_i1(Co29_C281),
            .Ck_j0(Co30_C290), .Ck_j1(Co30_C291), .Sk_01(S[31]), .Sk_i(N_220) );
sum_gen I176 ( .C_i(Co28_C270), .Cj_i0(Co29_C280), .Cj_i1(Co29_C281),
            .Ck_j0(Co30_C290), .Ck_j1(Co30_C291), .Sk_01(S[31]), .Sk_i(N_219) );
sum_gen I177 ( .C_i(C27_C231), .Cj_i0(Co28_C270), .Cj_i1(Co28_C271),
            .Ck_j0(Co29_C280), .Ck_j1(Co29_C281), .Sk_01(S[30]), .Sk_i(N_217) );
sum_gen I178 ( .C_i(C27_C230), .Cj_i0(Co28_C270), .Cj_i1(Co28_C271),
            .Ck_j0(Co29_C280), .Ck_j1(Co29_C281), .Sk_01(S[30]), .Sk_i(N_218) );
sum_gen I179 ( .C_i(gnd), .Cj_i0(C27_C231), .Cj_i1(gnd), .Ck_j0(Co28_C270),
            .Ck_j1(Co28_C271), .Sk_01(S[29]), .Sk_i(N_215) );
sum_gen I180 ( .C_i(gnd), .Cj_i0(C27_C230), .Cj_i1(gnd), .Ck_j0(Co28_C270),
            .Ck_j1(Co28_C271), .Sk_01(S[29]), .Sk_i(N_216) );
sum_gen I181 ( .C_i(Co20_C191), .Cj_i0(Co21_C200), .Cj_i1(Co21_C201),
            .Ck_j0(Co22_C210), .Ck_j1(Co22_C211), .Sk_01(S[23]), .Sk_i(N_225) );
sum_gen I182 ( .C_i(Co20_C190), .Cj_i0(Co21_C200), .Cj_i1(Co21_C201),
            .Ck_j0(Co22_C210), .Ck_j1(Co22_C211), .Sk_01(S[23]), .Sk_i(N_226) );
sum_gen I183 ( .C_i(C19_C151), .Cj_i0(Co20_C190), .Cj_i1(Co20_C191),
            .Ck_j0(Co21_C200), .Ck_j1(Co21_C201), .Sk_01(S[22]), .Sk_i(N_223) );
sum_gen I184 ( .C_i(C19_C150), .Cj_i0(Co20_C190), .Cj_i1(Co20_C191),
            .Ck_j0(Co21_C200), .Ck_j1(Co21_C201), .Sk_01(S[22]), .Sk_i(N_224) );
sum_gen I185 ( .C_i(Carry15), .Cj_i0(C19_C150), .Cj_i1(C19_C151),
            .Ck_j0(Co20_C190), .Ck_j1(Co20_C191), .Sk_01(S[21]),
            .Sk_i(Sumi[21]) );
sum_gen I186 ( .C_i(gnd), .Cj_i0(Carry15), .Cj_i1(gnd), .Ck_j0(C19_C150),
            .Ck_j1(C19_C151), .Sk_01(S[20]), .Sk_i(Sumi[20]) );
sum_gen I187 ( .C_i(Co24_C231), .Cj_i0(Co25_C240), .Cj_i1(Co25_C241),
            .Ck_j0(Co26_C250), .Ck_j1(Co26_C251), .Sk_01(S[27]), .Sk_i(N_231) );
sum_gen I188 ( .C_i(Co24_C230), .Cj_i0(Co25_C240), .Cj_i1(Co25_C241),
            .Ck_j0(Co26_C250), .Ck_j1(Co26_C251), .Sk_01(S[27]), .Sk_i(N_232) );
sum_gen I189 ( .C_i(gnd), .Cj_i0(Co24_C231), .Cj_i1(gnd), .Ck_j0(Co25_C240),
            .Ck_j1(Co25_C241), .Sk_01(S[26]), .Sk_i(N_229) );
sum_gen I190 ( .C_i(gnd), .Cj_i0(Co24_C230), .Cj_i1(gnd), .Ck_j0(Co25_C240),
            .Ck_j1(Co25_C241), .Sk_01(S[26]), .Sk_i(N_230) );
sum_gen I191 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Co24_C231),
            .Ck_j1(gnd), .Sk_01(S[25]), .Sk_i(N_227) );
sum_gen I192 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Co24_C230),
            .Ck_j1(gnd), .Sk_01(S[25]), .Sk_i(N_228) );
sum_gen I193 ( .C_i(Carry15), .Cj_i0(C19_C150), .Cj_i1(C19_C151),
            .Ck_j0(C23_C190), .Ck_j1(C23_C191), .Sk_01(S[24]),
            .Sk_i(Sumi[24]) );
sum_gen I194 ( .C_i(Co16_C151), .Cj_i0(Co17_C160), .Cj_i1(Co17_C161),
            .Ck_j0(Co18_C170), .Ck_j1(Co18_C171), .Sk_01(S[19]), .Sk_i(N_233) );
sum_gen I195 ( .C_i(Co16_C150), .Cj_i0(Co17_C160), .Cj_i1(Co17_C161),
            .Ck_j0(Co18_C170), .Ck_j1(Co18_C171), .Sk_01(S[19]), .Sk_i(N_234) );
sum_gen I196 ( .C_i(Carry15a), .Cj_i0(Co16_C150), .Cj_i1(Co16_C151),
            .Ck_j0(Co17_C160), .Ck_j1(Co17_C161), .Sk_01(S[18]),
            .Sk_i(Sumi[18]) );
sum_gen I197 ( .C_i(gnd), .Cj_i0(Carry15a), .Cj_i1(gnd), .Ck_j0(Co16_C150),
            .Ck_j1(Co16_C151), .Sk_01(S[17]), .Sk_i(Sumi[17]) );
sum_gen I198 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Carry15a), .Ck_j1(gnd),
            .Sk_01(S[16]), .Sk_i(Sumi[16]) );
sum_gen I149 ( .C_i(Co12_C111), .Cj_i0(Co13_C120), .Cj_i1(Co13_C121),
            .Ck_j0(Co14_C130), .Ck_j1(Co14_C131), .Sk_01(S[15]), .Sk_i(N_211) );
sum_gen I150 ( .C_i(Co12_C110), .Cj_i0(Co13_C120), .Cj_i1(Co13_C121),
            .Ck_j0(Co14_C130), .Ck_j1(Co14_C131), .Sk_01(S[15]), .Sk_i(N_212) );
sum_gen I151 ( .C_i(gnd), .Cj_i0(Co12_C111), .Cj_i1(gnd), .Ck_j0(Co13_C120),
            .Ck_j1(Co13_C121), .Sk_01(S[14]), .Sk_i(N_209) );
sum_gen I152 ( .C_i(gnd), .Cj_i0(Co12_C110), .Cj_i1(gnd), .Ck_j0(Co13_C120),
            .Ck_j1(Co13_C121), .Sk_01(S[14]), .Sk_i(N_210) );
sum_gen I153 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Co12_C111),
            .Ck_j1(gnd), .Sk_01(S[13]), .Sk_i(N_207) );
sum_gen I154 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Co12_C110),
            .Ck_j1(gnd), .Sk_01(S[13]), .Sk_i(N_208) );
sum_gen I155 ( .C_i(Carry3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
            .Ck_j1(C11_C71), .Sk_01(S[12]), .Sk_i(Sumi[12]) );
sum_gen I143 ( .C_i(Co8_C71), .Cj_i0(Co9_C80), .Cj_i1(Co9_C81), .Ck_j0(Co10_C90),
            .Ck_j1(Co10_C91), .Sk_01(S[11]), .Sk_i(N_201) );
sum_gen I144 ( .C_i(Co8_C70), .Cj_i0(Co9_C80), .Cj_i1(Co9_C81), .Ck_j0(Co10_C90),
            .Ck_j1(Co10_C91), .Sk_01(S[11]), .Sk_i(N_202) );
sum_gen I145 ( .C_i(gnd), .Cj_i0(Co8_C71), .Cj_i1(gnd), .Ck_j0(Co9_C80),
            .Ck_j1(Co9_C81), .Sk_01(S[10]), .Sk_i(N_204) );
sum_gen I146 ( .C_i(gnd), .Cj_i0(Co8_C70), .Cj_i1(gnd), .Ck_j0(Co9_C80),
            .Ck_j1(Co9_C81), .Sk_01(S[10]), .Sk_i(N_203) );
sum_gen I147 ( .C_i(Carry3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(Co8_C70),
            .Ck_j1(Co8_C71), .Sk_01(S[9]), .Sk_i(Sumi[9]) );
sum_gen I148 ( .C_i(gnd), .Cj_i0(Carry3a), .Cj_i1(gnd), .Ck_j0(C7_C30),
            .Ck_j1(C7_C31), .Sk_01(S[8]), .Sk_i(Sumi[8]) );
sum_gen I138 ( .C_i(Co4_C31), .Cj_i0(Co5_C40), .Cj_i1(Co5_C41), .Ck_j0(Co6_C50),
            .Ck_j1(Co6_C51), .Sk_01(S[7]), .Sk_i(N_206) );
sum_gen I139 ( .C_i(Co4_C30), .Cj_i0(Co5_C40), .Cj_i1(Co5_C41), .Ck_j0(Co6_C50),
            .Ck_j1(Co6_C51), .Sk_01(S[7]), .Sk_i(N_205) );
sum_gen I140 ( .C_i(Carry3), .Cj_i0(Co4_C30), .Cj_i1(Co4_C31), .Ck_j0(Co5_C40),
            .Ck_j1(Co5_C41), .Sk_01(S[6]), .Sk_i(Sumi[6]) );
sum_gen I141 ( .C_i(gnd), .Cj_i0(Carry3), .Cj_i1(gnd), .Ck_j0(Co4_C30),
            .Ck_j1(Co4_C31), .Sk_01(S[5]), .Sk_i(Sumi[5]) );
sum_gen I142 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Carry3), .Ck_j1(gnd),
            .Sk_01(S[4]), .Sk_i(Sumi[4]) );
sum_gen I135 ( .C_i(Carry_0), .Cj_i0(Co1_C00), .Cj_i1(Co1_C01), .Ck_j0(Co2_C10),
            .Ck_j1(Co2_C11), .Sk_01(S[3]), .Sk_i(Sumi[3]) );
sum_gen I136 ( .C_i(Cin), .Cj_i0(Co0_Ci0), .Cj_i1(Co0_Ci1), .Ck_j0(Co1_C00),
            .Ck_j1(Co1_C01), .Sk_01(S[2]), .Sk_i(Sumi[2]) );
sum_gen I137 ( .C_i(gnd), .Cj_i0(Cin), .Cj_i1(gnd), .Ck_j0(Co0_Ci0),
            .Ck_j1(Co0_Ci1), .Sk_01(S[1]), .Sk_i(Sumi[1]) );
sum0 I132 ( .A(a[0]), .B(b[0]), .Cin(Cin), .s0(Sumi[0]) );

endmodule // sum32

`endif

`ifdef sum16
`else
`define sum16
module sum16( a , b, C11_C70, C11_C71, C7_C30, C7_C31, Cin, Co0_Ci0, Co0_Ci1,
              Co10_C90, Co10_C91, Co12_C110, Co12_C111, Co13_C120, Co13_C121,
              Co14_C130, Co14_C131, Co1_C00, Co1_C01, Co2_C10, Co2_C11,
              Co3_C20, Co3_C21, Co4_C30, Co4_C31, Co5_C40, Co5_C41, Co6_C50,
              Co6_C51, Co8_C70, Co8_C71, Co9_C80, Co9_C81, S, Carry3, Sumi );
 input [0:0] a;
 input [0:0] b;
input C11_C70, C11_C71, C7_C30, C7_C31;
output Carry3;
input Cin, Co0_Ci0, Co0_Ci1, Co10_C90, Co10_C91, Co12_C110, Co12_C111,
Co13_C120, Co13_C121, Co14_C130, Co14_C131, Co1_C00, Co1_C01, Co2_C10,
Co2_C11, Co3_C20, Co3_C21, Co4_C30, Co4_C31, Co5_C40, Co5_C41, Co6_C50,
Co6_C51, Co8_C70, Co8_C71, Co9_C80, Co9_C81;
 input [15:0] S;
 output [15:0] Sumi;
wire Carry_0;
wire N_39;
wire N_40;
wire N_33;
wire N_34;
wire N_35;
wire N_36;
wire N_37;
wire N_38;
wire N_29;
wire N_30;
wire N_31;
wire N_32;
wire Carry3a;
supply0 gnd;

sum2_gen I107 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Carry3), .Ck_j1(gnd),
             .Sk_0(N_39), .Sk_1(N_40), .Sk_i(Sumi[7]) );
sum2_gen I108 ( .C_i(gnd), .Cj_i0(Carry3a), .Cj_i1(gnd), .Ck_j0(C7_C30),
             .Ck_j1(C7_C31), .Sk_0(N_30), .Sk_1(N_29), .Sk_i(Sumi[11]) );
sum2_gen I109 ( .C_i(gnd), .Cj_i0(Carry3a), .Cj_i1(gnd), .Ck_j0(C7_C30),
             .Ck_j1(C7_C31), .Sk_0(N_31), .Sk_1(N_32), .Sk_i(Sumi[10]) );
sum2_gen I94 ( .C_i(Carry3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
            .Ck_j1(C11_C71), .Sk_0(N_38), .Sk_1(N_33), .Sk_i(Sumi[13]) );
sum2_gen I95 ( .C_i(Carry3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
            .Ck_j1(C11_C71), .Sk_0(N_37), .Sk_1(N_35), .Sk_i(Sumi[14]) );
sum2_gen I96 ( .C_i(Carry3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
            .Ck_j1(C11_C71), .Sk_0(N_36), .Sk_1(N_34), .Sk_i(Sumi[15]) );
cary_gen I110 ( .C_i(Carry_0), .Cj_i0(Co1_C00), .Cj_i1(Co1_C01), .Ck_j0(Co2_C10),
             .Ck_j1(Co2_C11), .Cm_i(Carry3a), .Cm_k0(Co3_C20),
             .Cm_k1(Co3_C21) );
cary_gen I111 ( .C_i(Carry_0), .Cj_i0(Co1_C00), .Cj_i1(Co1_C01), .Ck_j0(Co2_C10),
             .Ck_j1(Co2_C11), .Cm_i(Carry3), .Cm_k0(Co3_C20), .Cm_k1(Co3_C21) );
carry0 I81 ( .A(a[0]), .B(b[0]), .Cin(Cin), .Cout(Carry_0) );
sum_gen I104 ( .C_i(gnd), .Cj_i0(Co12_C111), .Cj_i1(gnd), .Ck_j0(Co13_C120),
            .Ck_j1(Co13_C121), .Sk_01(S[14]), .Sk_i(N_35) );
sum_gen I97 ( .C_i(Co12_C111), .Cj_i0(Co13_C120), .Cj_i1(Co13_C121),
           .Ck_j0(Co14_C130), .Ck_j1(Co14_C131), .Sk_01(S[15]), .Sk_i(N_34) );
sum_gen I98 ( .C_i(Co12_C110), .Cj_i0(Co13_C120), .Cj_i1(Co13_C121),
           .Ck_j0(Co14_C130), .Ck_j1(Co14_C131), .Sk_01(S[15]), .Sk_i(N_36) );
sum_gen I99 ( .C_i(Co4_C31), .Cj_i0(Co5_C40), .Cj_i1(Co5_C41), .Ck_j0(Co6_C50),
           .Ck_j1(Co6_C51), .Sk_01(S[7]), .Sk_i(N_40) );
sum_gen I100 ( .C_i(Co4_C30), .Cj_i0(Co5_C40), .Cj_i1(Co5_C41), .Ck_j0(Co6_C50),
            .Ck_j1(Co6_C51), .Sk_01(S[7]), .Sk_i(N_39) );
sum_gen I101 ( .C_i(Carry3), .Cj_i0(Co4_C30), .Cj_i1(Co4_C31), .Ck_j0(Co5_C40),
            .Ck_j1(Co5_C41), .Sk_01(S[6]), .Sk_i(Sumi[6]) );
sum_gen I102 ( .C_i(gnd), .Cj_i0(Carry3), .Cj_i1(gnd), .Ck_j0(Co4_C30),
            .Ck_j1(Co4_C31), .Sk_01(S[5]), .Sk_i(Sumi[5]) );
sum_gen I103 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Carry3), .Ck_j1(gnd),
            .Sk_01(S[4]), .Sk_i(Sumi[4]) );
sum_gen I105 ( .C_i(gnd), .Cj_i0(Co12_C110), .Cj_i1(gnd), .Ck_j0(Co13_C120),
            .Ck_j1(Co13_C121), .Sk_01(S[14]), .Sk_i(N_37) );
sum_gen I106 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Co12_C111),
            .Ck_j1(gnd), .Sk_01(S[13]), .Sk_i(N_33) );
sum_gen I83 ( .C_i(Carry_0), .Cj_i0(Co1_C00), .Cj_i1(Co1_C01), .Ck_j0(Co2_C10),
           .Ck_j1(Co2_C11), .Sk_01(S[3]), .Sk_i(Sumi[3]) );
sum_gen I84 ( .C_i(Cin), .Cj_i0(Co0_Ci0), .Cj_i1(Co0_Ci1), .Ck_j0(Co1_C00),
           .Ck_j1(Co1_C01), .Sk_01(S[2]), .Sk_i(Sumi[2]) );
sum_gen I85 ( .C_i(gnd), .Cj_i0(Cin), .Cj_i1(gnd), .Ck_j0(Co0_Ci0),
           .Ck_j1(Co0_Ci1), .Sk_01(S[1]), .Sk_i(Sumi[1]) );
sum_gen I86 ( .C_i(gnd), .Cj_i0(gnd), .Cj_i1(gnd), .Ck_j0(Co12_C110), .Ck_j1(gnd),
           .Sk_01(S[13]), .Sk_i(N_38) );
sum_gen I87 ( .C_i(Carry3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
           .Ck_j1(C11_C71), .Sk_01(S[12]), .Sk_i(Sumi[12]) );
sum_gen I88 ( .C_i(Co8_C71), .Cj_i0(Co9_C80), .Cj_i1(Co9_C81), .Ck_j0(Co10_C90),
           .Ck_j1(Co10_C91), .Sk_01(S[11]), .Sk_i(N_29) );
sum_gen I89 ( .C_i(Co8_C70), .Cj_i0(Co9_C80), .Cj_i1(Co9_C81), .Ck_j0(Co10_C90),
           .Ck_j1(Co10_C91), .Sk_01(S[11]), .Sk_i(N_30) );
sum_gen I90 ( .C_i(gnd), .Cj_i0(Co8_C71), .Cj_i1(gnd), .Ck_j0(Co9_C80),
           .Ck_j1(Co9_C81), .Sk_01(S[10]), .Sk_i(N_32) );
sum_gen I91 ( .C_i(gnd), .Cj_i0(Co8_C70), .Cj_i1(gnd), .Ck_j0(Co9_C80),
           .Ck_j1(Co9_C81), .Sk_01(S[10]), .Sk_i(N_31) );
sum_gen I92 ( .C_i(Carry3a), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(Co8_C70),
           .Ck_j1(Co8_C71), .Sk_01(S[9]), .Sk_i(Sumi[9]) );
sum_gen I93 ( .C_i(gnd), .Cj_i0(Carry3a), .Cj_i1(gnd), .Ck_j0(C7_C30),
           .Ck_j1(C7_C31), .Sk_01(S[8]), .Sk_i(Sumi[8]) );
sum0 I82 ( .A(a[0]), .B(b[0]), .Cin(Cin), .s0(Sumi[0]) );

endmodule // sum16

`endif

`ifdef carry16
`else
`define carry16
module carry16( a , b, Carry3, C11_C70, C11_C71, C7_C30, C7_C31, Co, Co0_Ci0,
                Co0_Ci1, Co10_C90, Co10_C91, Co12_C110, Co12_C111, Co13_C120,
                Co13_C121, Co14_C130, Co14_C131, Co1_C00, Co1_C01, Co2_C10,
                Co2_C11, Co3_C20, Co3_C21, Co4_C30, Co4_C31, Co5_C40, Co5_C41,
                Co6_C50, Co6_C51, Co8_C70, Co8_C71, Co9_C80, Co9_C81, S );
 input [15:0] a;
 input [15:0] b;
output C11_C70, C11_C71, C7_C30, C7_C31;
input Carry3;
output Co, Co0_Ci0, Co0_Ci1, Co10_C90, Co10_C91, Co12_C110, Co12_C111,
Co13_C120, Co13_C121, Co14_C130, Co14_C131, Co1_C00, Co1_C01, Co2_C10,
Co2_C11, Co3_C20, Co3_C21, Co4_C30, Co4_C31, Co5_C40, Co5_C41, Co6_C50,
Co6_C51, Co8_C70, Co8_C71, Co9_C80, Co9_C81;
 output [15:0] S;
wire Co7_C60;
wire Co7_C61;
wire Co11_C100;
wire Co11_C101;
wire C15_C110;
wire C15_C111;
wire Co15_C140;
wire Co15_C141;

sum_c0 s0 ( .Ax(a[0]), .Bx(b[0]), .Co_Ci0(Co0_Ci0), .Co_Ci1(Co0_Ci1) );
cary_gen I46 ( .C_i(Co8_C71), .Cj_i0(Co9_C80), .Cj_i1(Co9_C81), .Ck_j0(Co10_C90),
            .Ck_j1(Co10_C91), .Cm_i(C11_C71), .Cm_k0(Co11_C100),
            .Cm_k1(Co11_C101) );
cary_gen I47 ( .C_i(Co8_C70), .Cj_i0(Co9_C80), .Cj_i1(Co9_C81), .Ck_j0(Co10_C90),
            .Ck_j1(Co10_C91), .Cm_i(C11_C70), .Cm_k0(Co11_C100),
            .Cm_k1(Co11_C101) );
cary_gen I41 ( .C_i(Carry3), .Cj_i0(C7_C30), .Cj_i1(C7_C31), .Ck_j0(C11_C70),
            .Ck_j1(C11_C71), .Cm_i(Co), .Cm_k0(C15_C110), .Cm_k1(C15_C111) );
cary_gen I42 ( .C_i(Co12_C111), .Cj_i0(Co13_C120), .Cj_i1(Co13_C121),
            .Ck_j0(Co14_C130), .Ck_j1(Co14_C131), .Cm_i(C15_C111),
            .Cm_k0(Co15_C140), .Cm_k1(Co15_C141) );
cary_gen I43 ( .C_i(Co12_C110), .Cj_i0(Co13_C120), .Cj_i1(Co13_C121),
            .Ck_j0(Co14_C130), .Ck_j1(Co14_C131), .Cm_i(C15_C110),
            .Cm_k0(Co15_C140), .Cm_k1(Co15_C141) );
cary_gen I44 ( .C_i(Co4_C31), .Cj_i0(Co5_C40), .Cj_i1(Co5_C41), .Ck_j0(Co6_C50),
            .Ck_j1(Co6_C51), .Cm_i(C7_C31), .Cm_k0(Co7_C60), .Cm_k1(Co7_C61) );
cary_gen I45 ( .C_i(Co4_C30), .Cj_i0(Co5_C40), .Cj_i1(Co5_C41), .Ck_j0(Co6_C50),
            .Ck_j1(Co6_C51), .Cm_i(C7_C30), .Cm_k0(Co7_C60), .Cm_k1(Co7_C61) );
sum_c s4 ( .Ax(a[4]), .Bx(b[4]), .Co_Ci0(Co4_C30), .Co_Ci1(Co4_C31),
        .Sub_Sum(S[4]) );
sum_c s15 ( .Ax(a[15]), .Bx(b[15]), .Co_Ci0(Co15_C140), .Co_Ci1(Co15_C141),
         .Sub_Sum(S[15]) );
sum_c s14 ( .Ax(a[14]), .Bx(b[14]), .Co_Ci0(Co14_C130), .Co_Ci1(Co14_C131),
         .Sub_Sum(S[14]) );
sum_c s12 ( .Ax(a[12]), .Bx(b[12]), .Co_Ci0(Co12_C110), .Co_Ci1(Co12_C111),
         .Sub_Sum(S[12]) );
sum_c s13 ( .Ax(a[13]), .Bx(b[13]), .Co_Ci0(Co13_C120), .Co_Ci1(Co13_C121),
         .Sub_Sum(S[13]) );
sum_c s11 ( .Ax(a[11]), .Bx(b[11]), .Co_Ci0(Co11_C100), .Co_Ci1(Co11_C101),
         .Sub_Sum(S[11]) );
sum_c s10 ( .Ax(a[10]), .Bx(b[10]), .Co_Ci0(Co10_C90), .Co_Ci1(Co10_C91),
         .Sub_Sum(S[10]) );
sum_c s8 ( .Ax(a[8]), .Bx(b[8]), .Co_Ci0(Co8_C70), .Co_Ci1(Co8_C71),
        .Sub_Sum(S[8]) );
sum_c s9 ( .Ax(a[9]), .Bx(b[9]), .Co_Ci0(Co9_C80), .Co_Ci1(Co9_C81),
        .Sub_Sum(S[9]) );
sum_c s7 ( .Ax(a[7]), .Bx(b[7]), .Co_Ci0(Co7_C60), .Co_Ci1(Co7_C61),
        .Sub_Sum(S[7]) );
sum_c s6 ( .Ax(a[6]), .Bx(b[6]), .Co_Ci0(Co6_C50), .Co_Ci1(Co6_C51),
        .Sub_Sum(S[6]) );
sum_c s5 ( .Ax(a[5]), .Bx(b[5]), .Co_Ci0(Co5_C40), .Co_Ci1(Co5_C41),
        .Sub_Sum(S[5]) );
sum_c s3 ( .Ax(a[3]), .Bx(b[3]), .Co_Ci0(Co3_C20), .Co_Ci1(Co3_C21),
        .Sub_Sum(S[3]) );
sum_c s2 ( .Ax(a[2]), .Bx(b[2]), .Co_Ci0(Co2_C10), .Co_Ci1(Co2_C11),
        .Sub_Sum(S[2]) );
sum_c s1 ( .Ax(a[1]), .Bx(b[1]), .Co_Ci0(Co1_C00), .Co_Ci1(Co1_C01),
        .Sub_Sum(S[1]) );

endmodule // carry16

`endif

`ifdef jknn_ff
`else
`define jknn_ff
module jknn_ff( CLK , CLR, J, KNN, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input J, KNN;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(GND), .QZ(Q) );
frag_m I_2 ( .B1(Q), .B2(GND), .C1(GND), .C2(VCC), .D1(VCC), .D2(GND), .E1(VCC),
          .E2(Q), .NS(N_3), .OS(N_2), .OZ(N_1) );
frag_f I_1 ( .F1(VCC), .F2(KNN), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_3) );
frag_a QL1 ( .A1(J), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // jknn_ff

`endif

`ifdef dladinv
`else
`define dladinv
module dladinv( DATA , G, Q, QNN );
input DATA, G;
output Q, QNN;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply0 GND;
supply1 VCC;

frag_m I_2 ( .B1(Q), .B2(GND), .C1(DATA), .C2(GND), .D1(QNN), .D2(GND), .E1(VCC),
          .E2(DATA), .NS(N_2), .NZ(QNN), .OS(N_1), .OZ(Q) );
frag_f I_1 ( .F1(G), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );
frag_a QL1 ( .A1(GND), .A2(VCC), .A3(GND), .A4(VCC), .A5(GND), .A6(VCC), .AZ(N_1) );

endmodule // dladinv

`endif

`ifdef s_r_ltch
`else
`define s_r_ltch
module s_r_ltch( R , S1, S2, Q, QN );
output Q, QN;
input R, S1, S2;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;

frag_a I_2 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_1) );
frag_f I_1 ( .F1(S1), .F2(GND), .F3(S2), .F4(GND), .F5(VCC), .F6(Q), .FZ(QN) );
frag_m QL1 ( .B1(GND), .B2(GND), .C1(GND), .C2(GND), .D1(R), .D2(GND), .E1(GND),
          .E2(VCC), .NS(QN), .NZ(Q), .OS(N_1) );

endmodule // s_r_ltch

`endif

`ifdef bank259
`else
`define bank259
module bank259( CLRNN , D0, D1, D2, D3, D4, D5, D6, D7, DATA, GNN, Q0, Q1, Q2, Q3,
                Q4, Q5, Q6, Q7 );
input CLRNN, D0, D1, D2, D3, D4, D5, D6, D7, DATA, GNN;
output Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7;

ltch259 I_1 ( .CLRNN(CLRNN), .DATA(DATA), .DECIN(D7), .GNN(GNN), .Q(Q7) );
ltch259 I_2 ( .CLRNN(CLRNN), .DATA(DATA), .DECIN(D6), .GNN(GNN), .Q(Q6) );
ltch259 I_3 ( .CLRNN(CLRNN), .DATA(DATA), .DECIN(D5), .GNN(GNN), .Q(Q5) );
ltch259 I_4 ( .CLRNN(CLRNN), .DATA(DATA), .DECIN(D4), .GNN(GNN), .Q(Q4) );
ltch259 I_5 ( .CLRNN(CLRNN), .DATA(DATA), .DECIN(D3), .GNN(GNN), .Q(Q3) );
ltch259 I_6 ( .CLRNN(CLRNN), .DATA(DATA), .DECIN(D2), .GNN(GNN), .Q(Q2) );
ltch259 I_7 ( .CLRNN(CLRNN), .DATA(DATA), .DECIN(D1), .GNN(GNN), .Q(Q1) );
ltch259 I_8 ( .CLRNN(CLRNN), .DATA(DATA), .DECIN(D0), .GNN(GNN), .Q(Q0) );

endmodule // bank259

`endif

`ifdef a169
`else
`define a169
module a169( QA , QB, UPDWN, A, ANN, OUTB );
output A, ANN, OUTB;
input QA, QB, UPDWN;
parameter ql_gate = `LOGIC;
supply0 GND;
supply1 VCC;

frag_m I_2 ( .B1(VCC), .B2(GND), .C1(GND), .C2(VCC), .D1(GND), .D2(VCC), .E1(GND),
          .E2(VCC), .NS(A), .OS(ANN), .OZ(OUTB) );
frag_f I_1 ( .F1(QA), .F2(GND), .F3(QB), .F4(GND), .F5(UPDWN), .F6(GND), .FZ(A) );
frag_a QL1 ( .A1(VCC), .A2(QA), .A3(VCC), .A4(QB), .A5(VCC), .A6(UPDWN), .AZ(ANN) );

endmodule // a169

`endif

`ifdef b169
`else
`define b169
module b169( A , ANN, QC, OUTC );
input A, ANN;
output OUTC;
input QC;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply0 GND;
supply1 VCC;

frag_m I_2 ( .B1(VCC), .B2(VCC), .C1(VCC), .C2(GND), .D1(VCC), .D2(ANN), .E1(VCC),
          .E2(A), .NS(N_1), .NZ(OUTC), .OS(N_2) );
frag_f I_1 ( .F1(VCC), .F2(GND), .F3(QC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_a QL1 ( .A1(VCC), .A2(VCC), .A3(VCC), .A4(VCC), .A5(VCC), .A6(VCC), .AZ(N_2) );

endmodule // b169

`endif

`ifdef rco169
`else
`define rco169
module rco169( A , ANN, ENT, QC, QD, RCO );
input A, ANN, ENT, QC, QD;
output RCO;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply0 GND;
supply1 VCC;

frag_m I_2 ( .B1(VCC), .B2(GND), .C1(GND), .C2(GND), .D1(GND), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .OS(N_2), .OZ(RCO) );
frag_f I_1 ( .F1(A), .F2(GND), .F3(QC), .F4(GND), .F5(QD), .F6(ENT), .FZ(N_1) );
frag_a QL1 ( .A1(ANN), .A2(QC), .A3(VCC), .A4(QD), .A5(VCC), .A6(ENT), .AZ(N_2) );

endmodule // rco169

`endif

`ifdef reg169
`else
`define reg169
module reg169( CLK , D_IN, DATA, EN, FDBK, LDNN, Q );
input CLK /* synthesis syn_isclock=1 */;
input D_IN, DATA, EN, FDBK, LDNN;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply0 GND;
supply1 VCC;
wire N_3;

frag_q QL1 ( .QC(CLK), .QD(N_1), .QR(GND), .QS(GND), .QZ(Q) );
frag_a I_2 ( .A1(LDNN), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );
frag_m I_1 ( .B1(DATA), .B2(GND), .C1(DATA), .C2(GND), .D1(FDBK), .D2(GND),
          .E1(VCC), .E2(FDBK), .NS(N_3), .OS(N_2), .OZ(N_1) );
frag_f QL2 ( .F1(VCC), .F2(D_IN), .F3(VCC), .F4(GND), .F5(EN), .F6(GND), .FZ(N_3) );

endmodule // reg169

`endif

`ifdef uplsbit
`else
`define uplsbit
module uplsbit( CLK , CLR, D, ENP, ENT, LOAD, Q0, Q1, Q2, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input D, ENP, ENT, LOAD;
output Q;
input Q0, Q1, Q2;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply0 GND;
supply1 VCC;

frag_f I_3 ( .F1(Q0), .F2(CLR), .F3(Q1), .F4(ENT), .F5(Q2), .F6(ENP), .FZ(N_3) );
frag_q I_2 ( .QC(CLK), .QD(N_1), .QR(GND), .QS(GND), .QZ(Q) );
frag_m I_1 ( .B1(Q), .B2(CLR), .C1(VCC), .C2(Q), .D1(D), .D2(GND), .E1(D), .E2(GND),
          .NS(N_3), .OS(N_2), .OZ(N_1) );
frag_a QL1 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(CLR), .A5(VCC), .A6(LOAD), .AZ(N_2) );

endmodule // uplsbit

`endif

`ifdef uplabit
`else
`define uplabit
module uplabit( CLK , CLR, D, ENP, ENT, LOAD, Q0, Q1, Q2, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input D, ENP, ENT, LOAD;
output Q;
input Q0, Q1, Q2;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(GND), .QZ(Q) );
frag_f I_2 ( .F1(Q0), .F2(ENP), .F3(Q1), .F4(ENT), .F5(Q2), .F6(GND), .FZ(N_3) );
frag_m I_1 ( .B1(Q), .B2(GND), .C1(VCC), .C2(Q), .D1(D), .D2(GND), .E1(D), .E2(GND),
          .NS(N_3), .OS(N_2), .OZ(N_1) );
frag_a QL1 ( .A1(VCC), .A2(LOAD), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // uplabit

`endif

`ifdef muxde2x0
`else
`define muxde2x0
module muxde2x0( A1 , A2, B1, B2, GNN, SEL, Y1, Y2 );
input A1, A2, B1, B2, GNN, SEL;
output Y1, Y2;
parameter ql_gate = `LOGIC;
supply0 GND;
supply1 VCC;
wire N_1;
wire N_2;

frag_f I_2 ( .F1(SEL), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );
frag_m I_1 ( .B1(A1), .B2(GNN), .C1(B1), .C2(GNN), .D1(A2), .D2(GNN), .E1(B2),
          .E2(GNN), .NS(N_2), .NZ(Y2), .OS(N_1), .OZ(Y1) );
frag_a QL1 ( .A1(GND), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_1) );

endmodule // muxde2x0

`endif

`ifdef mux4x0e
`else
`define mux4x0e
module mux4x0e( A , B, C, D, GNN, S0, S1, Q );
input A, B, C, D, GNN;
output Q;
input S0, S1;
parameter ql_gate = `LOGIC;
supply0 GND;
wire N_1;
wire N_2;
supply1 VCC;

frag_f I_2 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );
frag_m I_1 ( .B1(A), .B2(GNN), .C1(B), .C2(GNN), .D1(C), .D2(GNN), .E1(D), .E2(GNN),
          .NS(N_2), .OS(N_1), .OZ(Q) );
frag_a QL1 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_1) );

endmodule // mux4x0e

`endif

`ifdef t148a2
`else
`define t148a2
module t148a2( EI , P4, P5, P6, P7, A2 );
output A2;
input EI, P4, P5, P6, P7;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(GND), .QD(A2), .QR(GND), .QS(GND) );
frag_m I_2 ( .B1(GND), .B2(VCC), .C1(P4), .C2(GND), .D1(VCC), .D2(GND), .E1(VCC),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(A2) );
frag_f I_1 ( .F1(P5), .F2(GND), .F3(P6), .F4(GND), .F5(P7), .F6(GND), .FZ(N_1) );
frag_a QL1 ( .A1(EI), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // t148a2

`endif

`ifdef t148a1
`else
`define t148a1
module t148a1( EI , P2, P3, P4, P5, P6, P7, A1 );
output A1;
input EI, P2, P3, P4, P5, P6, P7;
wire N_1;
wire N_2;
wire N_3;

or4i0 QL1 ( .A(EI), .B(N_3), .C(N_2), .D(N_1), .Q(A1) );
and4i0 QL2 ( .A(P3), .B(P2), .C(P7), .D(P6), .Q(N_3) );
and3i1 QL3 ( .A(P7), .B(P6), .C(P4), .Q(N_2) );
and3i1 QL4 ( .A(P6), .B(P7), .C(P5), .Q(N_1) );

endmodule // t148a1

`endif

`ifdef t148ao
`else
`define t148ao
module t148ao( EI , P1, P2, P3, P4, P5, P6, P7, A0 );
output A0;
input EI, P1, P2, P3, P4, P5, P6, P7;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;

xor2i0 QL1 ( .A(N_2), .B(N_1), .Q(A0) );
or3i0 QL2 ( .A(N_5), .B(N_4), .C(N_3), .Q(N_1) );
and4i2 QL3 ( .A(N_2), .B(P6), .C(P5), .D(EI), .Q(N_3) );
and5i2 QL4 ( .A(N_2), .B(P4), .C(P6), .D(P3), .E(EI), .Q(N_4) );
and6i2 QL5 ( .A(N_2), .B(P2), .C(P4), .D(P6), .E(P1), .F(EI), .Q(N_5) );
or2i0 QL6 ( .A(EI), .B(P7), .Q(N_2) );

endmodule // t148ao

`endif

`ifdef t138f3
`else
`define t138f3
module t138f3( A , B, C, EN, ENOUT, Y1, Y5 );
input A, B, C, EN;
output ENOUT, Y1, Y5;
parameter ql_gate = `LOGIC;
wire N_1;
supply1 VCC;
supply0 GND;

frag_q I_3 ( .QC(GND), .QD(N_1), .QR(GND), .QS(VCC) );
frag_m I_2 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(VCC), .D2(EN), .E1(VCC),
          .E2(EN), .NS(Y5), .NZ(ENOUT), .OS(Y1), .OZ(N_1) );
frag_f I_1 ( .F1(A), .F2(B), .F3(VCC), .F4(EN), .F5(C), .F6(EN), .FZ(Y5) );
frag_a QL1 ( .A1(A), .A2(EN), .A3(VCC), .A4(B), .A5(VCC), .A6(C), .AZ(Y1) );

endmodule // t138f3

`endif

`ifdef t138f2
`else
`define t138f2
module t138f2( A , B, C, EN, Y0, Y3, Y6 );
input A, B, C, EN;
output Y0, Y3, Y6;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(GND), .QD(Y3), .QR(GND), .QS(GND) );
frag_m I_2 ( .B1(VCC), .B2(VCC), .C1(A), .C2(C), .D1(GND), .D2(VCC), .E1(C), .E2(A),
          .NS(N_1), .NZ(Y6), .OS(Y0), .OZ(Y3) );
frag_f I_1 ( .F1(B), .F2(GND), .F3(EN), .F4(GND), .F5(EN), .F6(GND), .FZ(N_1) );
frag_a QL1 ( .A1(EN), .A2(A), .A3(EN), .A4(B), .A5(EN), .A6(C), .AZ(Y0) );

endmodule // t138f2

`endif

`ifdef t138f1
`else
`define t138f1
module t138f1( A , B, C, EN, Y2, Y4, Y7 );
input A, B, C, EN;
output Y2, Y4, Y7;
parameter ql_gate = `LOGIC;
supply0 GND;
wire N_1;
supply1 VCC;

frag_m I_2 ( .B1(VCC), .B2(VCC), .C1(C), .C2(B), .D1(GND), .D2(VCC), .E1(B), .E2(C),
          .NS(N_1), .NZ(Y2), .OS(Y7), .OZ(Y4) );
frag_f I_1 ( .F1(VCC), .F2(A), .F3(VCC), .F4(GND), .F5(VCC), .F6(EN), .FZ(N_1) );
frag_a QL1 ( .A1(A), .A2(EN), .A3(B), .A4(GND), .A5(C), .A6(GND), .AZ(Y7) );

endmodule // t138f1

`endif

`ifdef dladc
`else
`define dladc
module dladc( C1NN , C2NN, CLR, D1, D2, Q1, Q2 );
input C1NN, C2NN, CLR, D1, D2;
output Q1, Q2;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply0 GND;
supply1 VCC;

frag_f I_2 ( .F1(VCC), .F2(C1NN), .F3(VCC), .F4(C2NN), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_m I_1 ( .B1(Q1), .B2(CLR), .C1(D1), .C2(CLR), .D1(Q2), .D2(CLR), .E1(D2),
          .E2(CLR), .NS(N_1), .NZ(Q2), .OS(N_2), .OZ(Q1) );
frag_a QL1 ( .A1(GND), .A2(VCC), .A3(GND), .A4(VCC), .A5(GND), .A6(VCC), .AZ(N_2) );

endmodule // dladc

`endif

`ifdef jknffpc
`else
`define jknffpc
module jknffpc( CLK , CLR, J, K, PRE, Q );
input CLK /* synthesis syn_isclock=1 */;
input CLR /* synthesis syn_isclock=1 */;
input PRE /* synthesis syn_isclock=1 */;
input J, K;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(PRE), .QZ(Q) );
frag_m I_2 ( .B1(Q), .B2(GND), .C1(GND), .C2(VCC), .D1(VCC), .D2(GND), .E1(VCC),
          .E2(Q), .NS(N_3), .OS(N_2), .OZ(N_1) );
frag_f I_1 ( .F1(VCC), .F2(K), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_3) );
frag_a QL1 ( .A1(J), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // jknffpc

`endif

`ifdef frag_q
`else
`define frag_q
module frag_q( QC , QD, QR, QS, QZ );
input QD, QC, QR, QS;
output QZ;
parameter ql_frag = 1;
 reg QZ;
`ifdef synthesis
 always @ (posedge QC or posedge QR or posedge QS) 
     if (QR)
        #1 QZ = 1'b0;
     else if (QS)
        #1 QZ = 1'b1;
     else #1 QZ = QD;
`else
  always @ (QR or QS) begin
      if (QR)
         #1 assign QZ = 1'b0;
      else if (QS)
         #1 assign QZ = 1'b1;
      else
         #1 deassign QZ;
  end
  always @ (posedge QC)
         QZ = #1 QD;
  initial begin
    #1;
    if (QR)
         #1 assign QZ = 1'b0;
    else if (QS)
         #1 assign QZ = 1'b1;
  end
 `endif

endmodule // frag_q

`endif

`ifdef frag_f
`else
`define frag_f
module frag_f( F1 , F2, F3, F4, F5, F6, FZ );
input F1, F2, F3, F4, F5, F6;
output FZ;
parameter ql_frag = 1;
 assign #1 FZ = F1 & ~F2 & F3 & ~F4 & F5 & ~F6;

endmodule // frag_f

`endif

`ifdef frag_m
`else
`define frag_m
module frag_m( B1 , B2, C1, C2, D1, D2, E1, E2, NS, OS, NZ, OZ );
input B1, B2, C1, C2, D1, D2, E1, E2, NS;
output NZ;
input OS;
output OZ;
parameter ql_frag = 1;
 assign #1 NZ = NS ? (E1 & ~E2):(D1 & ~D2);
 assign #1 OZ = OS ? NZ:(NS ? (C1 & ~C2):(B1 & ~B2));

endmodule // frag_m

`endif

`ifdef frag_a
`else
`define frag_a
module frag_a( A1 , A2, A3, A4, A5, A6, AZ );
input A1, A2, A3, A4, A5, A6;
output AZ;
parameter ql_frag = 1;
 assign #1 AZ = A1 & ~A2 & A3 & ~A4 & A5 & ~A6;

endmodule // frag_a

`endif

`ifdef tri_inv
`else
`define tri_inv
module tri_inv( IN1 , IN2, IN3, OUT1, OUT2, OUT3 );
input IN1, IN2, IN3;
output OUT1, OUT2, OUT3;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;

frag_f I_2 ( .F1(VCC), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(IN3), .FZ(OUT3) );
frag_m I_1 ( .B1(GND), .B2(VCC), .C1(GND), .C2(VCC), .D1(VCC), .D2(IN2), .E1(VCC),
          .E2(IN2), .NS(OUT3), .NZ(OUT2), .OS(OUT1) );
frag_a QL1 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(IN1), .AZ(OUT1) );

endmodule // tri_inv

`endif

`ifdef bicell2
`else
`define bicell2
module bicell2( I1 , I2, IC, IE, IQE, IR, IQ, IZ, IP );
input I1, I2, IC, IE;
inout IP;
output IQ;
input IQE, IR;
output IZ;
parameter syn_macro = 1;
parameter ql_frag = 1;
reg IQ;
 assign #1 IP = IE ? (~I1 | I2):1'bz;
 assign #1 IZ = IP;
`ifdef synthesis
  always @ (posedge IC or posedge IR) 
     if (IR)
        #1 IQ = 1'b0;
     else if (IQE) 
        #1 IQ = IP;
`else
  always @ (posedge IC)
     if (~IR & IQE)
        #1 IQ = IP;
  always @ (IR) 
    #1 IQ = 1'b0;
 `endif

endmodule // bicell2

`endif

`ifdef incell2
`else
`define incell2
module incell2( IC , IP, IQE, IR, IN, IQ, IZ );
input IC;
output IN;
input IP;
output IQ;
input IQE, IR;
output IZ;
parameter syn_macro = 1;
parameter ql_frag = 1;
reg IQ;
 assign #1 IN = ~IP;
 assign #1 IZ = IP;
`ifdef synthesis
  always @ (posedge IC or posedge IR) 
     if (IR)
        #1 IQ = 1'b0;
     else if (IQE) 
        #1 IQ = IP;
`else
  always @ (posedge IC)
     if (~IR & IQE)
        #1 IQ = IP;
  always @ (IR) 
    #1 IQ = 1'b0;
 `endif

endmodule // incell2

`endif

`ifdef bufcell
`else
`define bufcell
module bufcell( IC , IZ );
input IC;
output IZ;
parameter ql_frag = 1;
 assign #1 IZ = IC;

endmodule // bufcell

`endif

`ifdef ckcell2
`else
`define ckcell2
module ckcell2( IP , IQC, IQE, IR, IC, IN, IQ, IZ );
output IC, IN;
input IP;
output IQ;
input IQC, IQE, IR;
output IZ;
parameter syn_macro = 1;
parameter ql_frag = 1;
reg IQ;
 assign #1 IN = ~IP;
 assign #1 IZ = IP;
 assign #1 IC = IP;
`ifdef synthesis
  always @ (posedge IQC or posedge IR) 
     if (IR)
        #1 IQ = 1'b0;
     else if (IQE) 
        #1 IQ = IP;
`else
  always @ (posedge IQC)
     if (~IR & IQE)
        #1 IQ = IP;
  always @ (IR) 
    #1 IQ = 1'b0;
 `endif

endmodule // ckcell2

`endif

`ifdef shiftbit
`else
`define shiftbit
module shiftbit( CLK , CLR, D, EN, LOAD, SI, Q );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input D, EN, LOAD;
output Q;
input SI;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;
wire N_1;
wire N_2;
wire N_3;

frag_a I_3 ( .A1(LOAD), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_1) );
frag_f I_2 ( .F1(EN), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );
frag_m I_1 ( .B1(Q), .B2(GND), .C1(SI), .C2(GND), .D1(D), .D2(GND), .E1(D), .E2(GND),
          .NS(N_2), .OS(N_1), .OZ(N_3) );
frag_q QL1 ( .QC(CLK), .QD(N_3), .QR(CLR), .QS(GND), .QZ(Q) );

endmodule // shiftbit

`endif

`ifdef bishbit
`else
`define bishbit
module bishbit( CLK , CLR, D, LSI, RSI, S0, S1, Q );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input D, LSI;
output Q;
input RSI, S0, S1;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;
wire N_1;
wire N_2;
wire N_3;

frag_a I_3 ( .A1(S1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_1) );
frag_f I_2 ( .F1(S0), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );
frag_m I_1 ( .B1(Q), .B2(GND), .C1(RSI), .C2(GND), .D1(LSI), .D2(GND), .E1(D),
          .E2(GND), .NS(N_2), .OS(N_1), .OZ(N_3) );
frag_q QL1 ( .QC(CLK), .QD(N_3), .QR(CLR), .QS(GND), .QZ(Q) );

endmodule // bishbit

`endif

`ifdef bicell
`else
`define bicell
module bicell( I1 , I2, IE, IZ, IP );
input I1, I2, IE;
inout IP;
output IZ;
parameter ql_frag = 1;
 assign #1 IP = IE ? (~I1 | I2):1'bz;
 assign #1 IZ = IP;

endmodule // bicell

`endif

`ifdef incell
`else
`define incell
module incell( IP , IN, IZ );
output IN;
input IP;
output IZ;
parameter ql_frag = 1;
 assign #1 IN = ~IP;
 assign #1 IZ = IP;

endmodule // incell

`endif

`ifdef ckcell
`else
`define ckcell
module ckcell( IP , IC, IN, IZ );
output IC, IN;
input IP;
output IZ;
parameter ql_frag = 1;
 assign #1 IN = ~IP;
 assign #1 IZ = IP;
 assign #1 IC = IP;

endmodule // ckcell

`endif

`ifdef udcnt3b
`else
`define udcnt3b
module udcnt3b( CLK , CLR, ENP, ENT, UP, Q, RCO );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input ENP, ENT;
 output [0:2] Q;
output RCO;
input UP;
supply1 VCC;
supply0 GND;

updnbitb QL4 ( .CLK(CLK), .CLR(CLR), .D0(GND), .D1(GND), .ENP(ENP), .ENT(ENT),
            .Q(Q[0]), .U0(VCC), .U1(VCC), .UP(UP) );
updnbitb QL3 ( .CLK(CLK), .CLR(CLR), .D0(Q[0]), .D1(GND), .ENP(ENP), .ENT(ENT),
            .Q(Q[1]), .U0(Q[0]), .U1(VCC), .UP(UP) );
updnbitb QL2 ( .CLK(CLK), .CLR(CLR), .D0(Q[0]), .D1(Q[1]), .ENP(ENP), .ENT(ENT),
            .Q(Q[2]), .U0(Q[0]), .U1(Q[1]), .UP(UP) );
updncarb QL1 ( .CO(RCO), .ENT(ENT), .Q0(Q[2]), .Q1(Q[1]), .Q2(Q[0]), .UP(UP) );

endmodule // udcnt3b

`endif

`ifdef udcnt3a
`else
`define udcnt3a
module udcnt3a( CLK , CLR, ENP, ENT, UP, Q, RCO );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input ENP, ENT;
 output [0:2] Q;
output RCO;
input UP;
supply1 VCC;
supply0 GND;

updnbita QL4 ( .CLK(CLK), .CLR(CLR), .D0(Q[0]), .D1(Q[1]), .ENP(ENP), .ENT(ENT),
            .Q(Q[2]), .U0(Q[0]), .U1(Q[1]), .UP(UP) );
updnbita QL3 ( .CLK(CLK), .CLR(CLR), .D0(Q[0]), .D1(GND), .ENP(ENP), .ENT(ENT),
            .Q(Q[1]), .U0(Q[0]), .U1(VCC), .UP(UP) );
updnbita QL2 ( .CLK(CLK), .CLR(CLR), .D0(GND), .D1(GND), .ENP(ENP), .ENT(ENT),
            .Q(Q[0]), .U0(VCC), .U1(VCC), .UP(UP) );
updncara QL1 ( .CO(RCO), .ENT(ENT), .Q0(Q[2]), .Q1(Q[1]), .Q2(Q[0]), .UP(UP) );

endmodule // udcnt3a

`endif

`ifdef uctxcar1
`else
`define uctxcar1
module uctxcar1( CLK , CLR, D, ENG, LOAD, Q, ACO1 );
output ACO1;
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [0:1] D;
input ENG, LOAD;
 input [0:1] Q;
wire N_1;
wire N_2;
wire N_3;

mux4x7 QL4 ( .A(N_2), .B(N_2), .C(N_3), .D(ACO1), .Q(N_1), .S0(ENG), .S1(LOAD) );
and2i1 QL3 ( .A(Q[1]), .B(Q[0]), .Q(N_3) );
and2i0 QL2 ( .A(D[0]), .B(D[1]), .Q(N_2) );
dffp QL1 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO1) );

endmodule // uctxcar1

`endif

`ifdef ucntx4c
`else
`define ucntx4c
module ucntx4c( CLK , CLR, D, ENG, ENP, ENT, LOAD, Q );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [0:3] D;
input ENG, ENP, ENT, LOAD;
 output [0:3] Q;
supply1 VCC;

upfxbit QL1 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
upfxbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(VCC) );
upfxbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[1]), .Q0(Q[0]), .Q1(VCC), .Q2(VCC) );
upfxbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[0]), .Q0(VCC), .Q1(VCC), .Q2(VCC) );

endmodule // ucntx4c

`endif

`ifdef ucntx4a
`else
`define ucntx4a
module ucntx4a( CLK , CLR, D, ENG, LOAD, Q, RCO );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [0:3] D;
input ENG, LOAD;
 output [0:3] Q;
output RCO;
supply0 GND;
supply1 VCC;

nand2i0 QL1 ( .A(Q[2]), .B(Q[3]), .Q(RCO) );
upfxbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENG(ENG), .ENP(GND), .ENT(GND),
           .LOAD(LOAD), .Q(Q[0]), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
upfxbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENG(ENG), .ENP(GND), .ENT(GND),
           .LOAD(LOAD), .Q(Q[1]), .Q0(Q[0]), .Q1(VCC), .Q2(VCC) );
upfxbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENG(ENG), .ENP(GND), .ENT(GND),
           .LOAD(LOAD), .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(VCC) );
upfxbit QL5 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENG(ENG), .ENP(GND), .ENT(GND),
           .LOAD(LOAD), .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );

endmodule // ucntx4a

`endif

`ifdef ucntx4b
`else
`define ucntx4b
module ucntx4b( CLK , CLR, D, ENG, ENP, ENT, LOAD, Q, RCO );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [0:3] D;
input ENG, ENP, ENT, LOAD;
 output [0:3] Q;
output RCO;
supply1 VCC;

nand5i1 QL1 ( .A(Q[0]), .B(Q[1]), .C(Q[2]), .D(Q[3]), .E(ENT), .Q(RCO) );
upfxbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
upfxbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(VCC) );
upfxbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[1]), .Q0(Q[0]), .Q1(VCC), .Q2(VCC) );
upfxbit QL5 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[0]), .Q0(VCC), .Q1(VCC), .Q2(VCC) );

endmodule // ucntx4b

`endif

`ifdef uctxcar2
`else
`define uctxcar2
module uctxcar2( CLK , CLR, D, ENG, LOAD, ACO1, ACO2 );
output ACO1, ACO2;
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [0:1] D;
input ENG, LOAD;
supply0 GND;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
supply1 VCC;

mux4x7 QL8 ( .A(N_4), .B(N_4), .C(N_5), .D(ACO2), .Q(N_1), .S0(ENG), .S1(LOAD) );
mux4x7 QL7 ( .A(N_4), .B(N_4), .C(N_5), .D(ACO1), .Q(N_2), .S0(ENG), .S1(LOAD) );
upfxbit QL6 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENG(ENG), .ENP(GND), .ENT(GND),
           .LOAD(LOAD), .Q(N_3), .Q0(N_6), .Q1(VCC), .Q2(VCC) );
upfxbit QL5 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENG(ENG), .ENP(GND), .ENT(GND),
           .LOAD(LOAD), .Q(N_6), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
and2i1 QL4 ( .A(N_3), .B(N_6), .Q(N_5) );
and2i0 QL3 ( .A(D[0]), .B(D[1]), .Q(N_4) );
dffp QL2 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO2) );
dffp QL1 ( .CLK(CLK), .D(N_2), .PRE(CLR), .Q(ACO1) );

endmodule // uctxcar2

`endif

`ifdef uctxcar3
`else
`define uctxcar3
module uctxcar3( CLK , CLR, D, ENG, LOAD, Q, ACO1, ACO2, ACO3 );
output ACO1, ACO2, ACO3;
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [0:1] D;
input ENG, LOAD;
 input [0:1] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;

mux4x7 QL8 ( .A(N_4), .B(N_4), .C(N_5), .D(ACO3), .Q(N_1), .S0(ENG), .S1(LOAD) );
mux4x7 QL7 ( .A(N_4), .B(N_4), .C(N_5), .D(ACO2), .Q(N_2), .S0(ENG), .S1(LOAD) );
mux4x7 QL6 ( .A(N_4), .B(N_4), .C(N_5), .D(ACO1), .Q(N_3), .S0(ENG), .S1(LOAD) );
and2i1 QL5 ( .A(Q[1]), .B(Q[0]), .Q(N_5) );
and2i0 QL4 ( .A(D[0]), .B(D[1]), .Q(N_4) );
dffp QL3 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO3) );
dffp QL2 ( .CLK(CLK), .D(N_2), .PRE(CLR), .Q(ACO2) );
dffp QL1 ( .CLK(CLK), .D(N_3), .PRE(CLR), .Q(ACO1) );

endmodule // uctxcar3

`endif

`ifdef uctlcar1
`else
`define uctlcar1
module uctlcar1( CLK , CLR, D, LOAD, Q, ACO1 );
output ACO1;
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [0:3] D;
input LOAD;
 input [0:3] Q;
supply0 GND;
supply1 VCC;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;

mux4x6 QL6 ( .A(VCC), .B(Q[3]), .C(D[3]), .D(VCC), .Q(N_1), .S0(N_4), .S1(N_5) );
and4i1 QL5 ( .A(LOAD), .B(N_3), .C(Q[2]), .D(N_2), .Q(N_4) );
and4i1 QL4 ( .A(D[0]), .B(D[1]), .C(D[2]), .D(LOAD), .Q(N_5) );
upflbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(N_3), .Q0(N_2), .Q1(VCC), .Q2(VCC) );
upflbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(N_2), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
dffp QL1 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO1) );

endmodule // uctlcar1

`endif

`ifdef ucntl4c
`else
`define ucntl4c
module ucntl4c( CLK , CLR, D, ENP, ENT, LOAD, Q );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [0:3] D;
input ENP, ENT, LOAD;
 output [0:3] Q;
supply1 VCC;

upflbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[0]), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
upflbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[1]), .Q0(Q[0]), .Q1(VCC), .Q2(VCC) );
upflbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(VCC) );
upflbit QL1 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );

endmodule // ucntl4c

`endif

`ifdef uctlcar3
`else
`define uctlcar3
module uctlcar3( CLK , CLR, D, LOAD, ACO1, ACO2, ACO3 );
output ACO1, ACO2, ACO3;
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [0:1] D;
input LOAD;
supply1 VCC;
supply0 GND;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;

and3i1 QL14 ( .A(D[0]), .B(D[1]), .C(LOAD), .Q(N_9) );
and3i1 QL13 ( .A(LOAD), .B(N_5), .C(N_4), .Q(N_6) );
and3i1 QL12 ( .A(D[0]), .B(D[1]), .C(LOAD), .Q(N_10) );
and3i1 QL11 ( .A(LOAD), .B(N_5), .C(N_4), .Q(N_7) );
and3i1 QL10 ( .A(LOAD), .B(N_5), .C(N_4), .Q(N_8) );
and3i1 QL9 ( .A(D[0]), .B(D[1]), .C(LOAD), .Q(N_11) );
mux4x0 QL8 ( .A(VCC), .B(GND), .C(GND), .D(VCC), .Q(N_1), .S0(N_6), .S1(N_9) );
mux4x0 QL7 ( .A(VCC), .B(GND), .C(GND), .D(VCC), .Q(N_2), .S0(N_7), .S1(N_10) );
mux4x0 QL6 ( .A(VCC), .B(GND), .C(GND), .D(VCC), .Q(N_3), .S0(N_8), .S1(N_11) );
upflbit QL5 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(N_5), .Q0(N_4), .Q1(VCC), .Q2(VCC) );
upflbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(N_4), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
dffp QL3 ( .CLK(CLK), .D(N_3), .PRE(CLR), .Q(ACO3) );
dffp QL2 ( .CLK(CLK), .D(N_2), .PRE(CLR), .Q(ACO2) );
dffp QL1 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO1) );

endmodule // uctlcar3

`endif

`ifdef uctlcar2
`else
`define uctlcar2
module uctlcar2( CLK , CLR, D, LOAD, ACO1, ACO2 );
output ACO1, ACO2;
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [0:1] D;
input LOAD;
supply0 GND;
supply1 VCC;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;

and3i1 QL10 ( .A(D[0]), .B(D[1]), .C(LOAD), .Q(N_7) );
and3i1 QL9 ( .A(LOAD), .B(N_4), .C(N_3), .Q(N_5) );
and3i1 QL8 ( .A(D[0]), .B(D[1]), .C(LOAD), .Q(N_8) );
and3i1 QL7 ( .A(LOAD), .B(N_4), .C(N_3), .Q(N_6) );
mux4x0 QL6 ( .A(VCC), .B(GND), .C(GND), .D(VCC), .Q(N_1), .S0(N_5), .S1(N_7) );
mux4x0 QL5 ( .A(VCC), .B(GND), .C(GND), .D(VCC), .Q(N_2), .S0(N_6), .S1(N_8) );
upflbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(N_4), .Q0(N_3), .Q1(VCC), .Q2(VCC) );
upflbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(N_3), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
dffp QL2 ( .CLK(CLK), .D(N_2), .PRE(CLR), .Q(ACO2) );
dffp QL1 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO1) );

endmodule // uctlcar2

`endif

`ifdef ucntl4b
`else
`define ucntl4b
module ucntl4b( CLK , CLR, D, ENP, ENT, LOAD, Q, RCO );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [0:3] D;
input ENP, ENT, LOAD;
 output [0:3] Q;
output RCO;
supply1 VCC;

upflbit QL5 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[0]), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
upflbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[1]), .Q0(Q[0]), .Q1(VCC), .Q2(VCC) );
upflbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(VCC) );
upflbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
nand5i1 QL1 ( .A(Q[0]), .B(Q[1]), .C(Q[2]), .D(Q[3]), .E(ENT), .Q(RCO) );

endmodule // ucntl4b

`endif

`ifdef ucntl4a
`else
`define ucntl4a
module ucntl4a( CLK , CLR, D, LOAD, Q, RCO );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [0:3] D;
input LOAD;
 output [0:3] Q;
output RCO;
supply0 GND;
supply1 VCC;

upflbit QL5 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(Q[0]), .Q0(VCC), .Q1(VCC), .Q2(VCC) );
upflbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(Q[1]), .Q0(Q[0]), .Q1(VCC), .Q2(VCC) );
upflbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(VCC) );
upflbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENP(GND), .ENT(GND), .LOAD(LOAD),
           .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
nand2i0 QL1 ( .A(Q[2]), .B(Q[3]), .Q(RCO) );

endmodule // ucntl4a

`endif

`ifdef uctecar1
`else
`define uctecar1
module uctecar1( CLK , CLR, ENG, Q, ACO1 );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
output ACO1;
input  ENG;
 input [0:3] Q;
wire N_1;
wire N_2;
supply0 GND;
wire N_3;
wire N_4;
supply1 VCC;

mux4x8 QL5 ( .A(VCC), .B(N_3), .C(VCC), .D(N_3), .Q(N_1), .S0(N_2), .S1(ENG) );
and3i0 QL4 ( .A(N_4), .B(Q[2]), .C(Q[3]), .Q(N_2) );
dffp QL3 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO1) );
upfebit QL2 ( .CLK(CLK), .CLR(CLR), .ENG(GND), .ENP(ENG), .ENT(GND), .Q(N_3),
           .Q0(VCC), .Q1(VCC), .Q2(VCC) );
upfebit QL1 ( .CLK(CLK), .CLR(CLR), .ENG(GND), .ENP(ENG), .ENT(GND), .Q(N_4),
           .Q0(N_3), .Q1(VCC), .Q2(VCC) );

endmodule // uctecar1

`endif

`ifdef ucnte4c
`else
`define ucnte4c
module ucnte4c( CLK , CLR, ENG, ENP, ENT, Q );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input ENG, ENP, ENT;
 output [0:3] Q;
supply1 VCC;

upfebit QL4 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(ENP), .ENT(ENT), .Q(Q[0]),
           .Q0(VCC), .Q1(VCC), .Q2(VCC) );
upfebit QL3 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(ENP), .ENT(ENT), .Q(Q[1]),
           .Q0(Q[0]), .Q1(VCC), .Q2(VCC) );
upfebit QL2 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(ENP), .ENT(ENT), .Q(Q[2]),
           .Q0(Q[0]), .Q1(Q[1]), .Q2(VCC) );
upfebit QL1 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(ENP), .ENT(ENT), .Q(Q[3]),
           .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );

endmodule // ucnte4c

`endif

`ifdef ucnte4b
`else
`define ucnte4b
module ucnte4b( CLK , CLR, ENG, ENP, ENT, Q, RCO );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input ENG, ENP, ENT;
 output [0:3] Q;
output RCO;
supply1 VCC;

upfebit QL5 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(ENP), .ENT(ENT), .Q(Q[0]),
           .Q0(VCC), .Q1(VCC), .Q2(VCC) );
upfebit QL4 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(ENP), .ENT(ENT), .Q(Q[1]),
           .Q0(Q[0]), .Q1(VCC), .Q2(VCC) );
upfebit QL3 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(ENP), .ENT(ENT), .Q(Q[2]),
           .Q0(Q[0]), .Q1(Q[1]), .Q2(VCC) );
upfebit QL2 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(ENP), .ENT(ENT), .Q(Q[3]),
           .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
nand5i1 QL1 ( .A(Q[0]), .B(Q[1]), .C(Q[2]), .D(Q[3]), .E(ENT), .Q(RCO) );

endmodule // ucnte4b

`endif

`ifdef ucnte4a
`else
`define ucnte4a
module ucnte4a( CLK , CLR, ENG, Q, RCO );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input ENG;
 output [0:3] Q;
output RCO;
supply1 VCC;
supply0 GND;

upfebit QL5 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(GND), .ENT(GND), .Q(Q[0]),
           .Q0(VCC), .Q1(VCC), .Q2(VCC) );
upfebit QL4 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(GND), .ENT(GND), .Q(Q[1]),
           .Q0(Q[0]), .Q1(VCC), .Q2(VCC) );
upfebit QL3 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(GND), .ENT(GND), .Q(Q[2]),
           .Q0(Q[0]), .Q1(Q[1]), .Q2(VCC) );
upfebit QL2 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(GND), .ENT(GND), .Q(Q[3]),
           .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
nand2i0 QL1 ( .A(Q[2]), .B(Q[3]), .Q(RCO) );

endmodule // ucnte4a

`endif

`ifdef upfecar2
`else
`define upfecar2
module upfecar2( CLK , CLR, ENG, ACO1, ACO2 );
output ACO1, ACO2;
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input ENG;
supply0 GND;
supply1 VCC;
wire N_1;
wire N_2;
wire N_3;
wire N_4;

mux4x8 QL6 ( .A(VCC), .B(N_3), .C(VCC), .D(N_3), .Q(N_2), .S0(N_4), .S1(ENG) );
mux4x8 QL5 ( .A(VCC), .B(N_3), .C(VCC), .D(N_3), .Q(N_1), .S0(N_4), .S1(ENG) );
dffp QL4 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO1) );
dffp QL3 ( .CLK(CLK), .D(N_2), .PRE(CLR), .Q(ACO2) );
upfebit QL2 ( .CLK(CLK), .CLR(CLR), .ENG(GND), .ENP(ENG), .ENT(GND), .Q(N_3),
           .Q0(VCC), .Q1(VCC), .Q2(VCC) );
upfebit QL1 ( .CLK(CLK), .CLR(CLR), .ENG(GND), .ENP(ENG), .ENT(GND), .Q(N_4),
           .Q0(N_3), .Q1(VCC), .Q2(VCC) );

endmodule // upfecar2

`endif

`ifdef upfecar3
`else
`define upfecar3
module upfecar3( CLK , CLR, ENG, ACO1, ACO2, ACO3 );
output ACO1, ACO2, ACO3;
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input ENG;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
supply0 GND;
supply1 VCC;

upfebit QL1 ( .CLK(CLK), .CLR(CLR), .ENG(GND), .ENP(ENG), .ENT(GND), .Q(N_1),
           .Q0(N_2), .Q1(VCC), .Q2(VCC) );
upfebit QL2 ( .CLK(CLK), .CLR(CLR), .ENG(GND), .ENP(ENG), .ENT(GND), .Q(N_2),
           .Q0(VCC), .Q1(VCC), .Q2(VCC) );
dffp QL3 ( .CLK(CLK), .D(N_4), .PRE(CLR), .Q(ACO2) );
dffp QL4 ( .CLK(CLK), .D(N_5), .PRE(CLR), .Q(ACO1) );
dffp QL5 ( .CLK(CLK), .D(N_3), .PRE(CLR), .Q(ACO3) );
mux4x8 QL6 ( .A(VCC), .B(N_2), .C(VCC), .D(N_2), .Q(N_5), .S0(N_1), .S1(ENG) );
mux4x8 QL7 ( .A(VCC), .B(N_2), .C(VCC), .D(N_2), .Q(N_4), .S0(N_1), .S1(ENG) );
mux4x8 QL8 ( .A(VCC), .B(N_2), .C(VCC), .D(N_2), .Q(N_3), .S0(N_1), .S1(ENG) );

endmodule // upfecar3

`endif

`ifdef ripbit
`else
`define ripbit
module ripbit( CI , CLK, CLR, CX, D, LOAD, CO, Q );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input CI;
output CO;
input CX, D, LOAD;
output Q;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(GND), .QZ(Q) );
frag_m I_2 ( .B1(Q), .B2(GND), .C1(VCC), .C2(Q), .D1(D), .D2(GND), .E1(D), .E2(GND),
          .NS(CO), .OS(N_2), .OZ(N_1) );
frag_f I_1 ( .F1(CI), .F2(GND), .F3(CX), .F4(GND), .F5(VCC), .F6(GND), .FZ(CO) );
frag_a QL1 ( .A1(LOAD), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // ripbit

`endif

`ifdef dctxcar1
`else
`define dctxcar1
module dctxcar1( CLK , CLR, D, ENG, LOAD, Q, ACO1 );
output ACO1;
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [1:0] D;
input ENG, LOAD;
 input [1:0] Q;
wire N_1;
wire N_2;
wire N_3;

dffp QL4 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO1) );
mux4x0 QL3 ( .A(ACO1), .B(N_3), .C(N_2), .D(N_2), .Q(N_1), .S0(ENG), .S1(LOAD) );
and2i2 QL2 ( .A(D[0]), .B(D[1]), .Q(N_2) );
and2i1 QL1 ( .A(Q[0]), .B(Q[1]), .Q(N_3) );

endmodule // dctxcar1

`endif

`ifdef dcntx4a
`else
`define dcntx4a
module dcntx4a( CLK , CLR, D, ENG, LOAD, Q, RCO );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [3:0] D;
input ENG, LOAD;
 output [3:0] Q;
output RCO;
supply1 VCC;
supply0 GND;

and2i2 QL5 ( .A(Q[2]), .B(Q[3]), .Q(RCO) );
dnfxbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENG(ENG), .ENP(VCC), .ENT(VCC),
           .LOAD(LOAD), .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
dnfxbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENG(ENG), .ENP(VCC), .ENT(VCC),
           .LOAD(LOAD), .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(GND) );
dnfxbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENG(ENG), .ENP(VCC), .ENT(VCC),
           .LOAD(LOAD), .Q(Q[1]), .Q0(Q[0]), .Q1(GND), .Q2(GND) );
dnfxbit QL1 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENG(ENG), .ENP(VCC), .ENT(VCC),
           .LOAD(LOAD), .Q(Q[0]), .Q0(GND), .Q1(GND), .Q2(GND) );

endmodule // dcntx4a

`endif

`ifdef dcntx4c
`else
`define dcntx4c
module dcntx4c( CLK , CLR, D, ENG, ENP, ENT, LOAD, Q );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [3:0] D;
input ENG, ENP, ENT, LOAD;
 output [3:0] Q;
supply0 GND;

dnfxbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
dnfxbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(GND) );
dnfxbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[1]), .Q0(Q[0]), .Q1(GND), .Q2(GND) );
dnfxbit QL1 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[0]), .Q0(GND), .Q1(GND), .Q2(GND) );

endmodule // dcntx4c

`endif

`ifdef dctxcar2
`else
`define dctxcar2
module dctxcar2( CLK , CLR, D, ENG, LOAD, ACO1, ACO2 );
output ACO1, ACO2;
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [1:0] D;
input ENG, LOAD;
wire N_1;
supply0 GND;
supply1 VCC;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;

dffp QL8 ( .CLK(CLK), .D(N_2), .PRE(CLR), .Q(ACO2) );
dffp QL7 ( .CLK(CLK), .D(N_3), .PRE(CLR), .Q(ACO1) );
and2i2 QL6 ( .A(D[0]), .B(D[1]), .Q(N_5) );
mux4x0 QL5 ( .A(ACO2), .B(N_1), .C(N_5), .D(N_5), .Q(N_2), .S0(ENG), .S1(LOAD) );
mux4x0 QL4 ( .A(ACO1), .B(N_1), .C(N_5), .D(N_5), .Q(N_3), .S0(ENG), .S1(LOAD) );
dnfxbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENG(ENG), .ENP(VCC), .ENT(VCC),
           .LOAD(LOAD), .Q(N_6), .Q0(GND), .Q1(GND), .Q2(GND) );
dnfxbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENG(ENG), .ENP(VCC), .ENT(VCC),
           .LOAD(LOAD), .Q(N_4), .Q0(N_6), .Q1(GND), .Q2(GND) );
and2i1 QL1 ( .A(N_6), .B(N_4), .Q(N_1) );

endmodule // dctxcar2

`endif

`ifdef dctxcar3
`else
`define dctxcar3
module dctxcar3( CLK , CLR, D, ENG, LOAD, Q, ACO1, ACO2, ACO3 );
output ACO1, ACO2, ACO3;
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [1:0] D;
input ENG, LOAD;
 input [1:0] Q;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;

dffp QL8 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO3) );
dffp QL7 ( .CLK(CLK), .D(N_2), .PRE(CLR), .Q(ACO2) );
dffp QL6 ( .CLK(CLK), .D(N_3), .PRE(CLR), .Q(ACO1) );
mux4x0 QL5 ( .A(ACO3), .B(N_5), .C(N_4), .D(N_4), .Q(N_1), .S0(ENG), .S1(LOAD) );
mux4x0 QL4 ( .A(ACO2), .B(N_5), .C(N_4), .D(N_4), .Q(N_2), .S0(ENG), .S1(LOAD) );
mux4x0 QL3 ( .A(ACO1), .B(N_5), .C(N_4), .D(N_4), .Q(N_3), .S0(ENG), .S1(LOAD) );
and2i2 QL2 ( .A(D[0]), .B(D[1]), .Q(N_4) );
and2i1 QL1 ( .A(Q[0]), .B(Q[1]), .Q(N_5) );

endmodule // dctxcar3

`endif

`ifdef dcntx4b
`else
`define dcntx4b
module dcntx4b( CLK , CLR, D, ENG, ENP, ENT, LOAD, Q, RCO );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [3:0] D;
input ENG, ENP, ENT, LOAD;
 output [3:0] Q;
output RCO;
supply0 GND;

and5i4 QL5 ( .A(ENT), .B(Q[0]), .C(Q[1]), .D(Q[2]), .E(Q[3]), .Q(RCO) );
dnfxbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
dnfxbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(GND) );
dnfxbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[1]), .Q0(Q[0]), .Q1(GND), .Q2(GND) );
dnfxbit QL1 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENG(ENG), .ENP(ENP), .ENT(ENT),
           .LOAD(LOAD), .Q(Q[0]), .Q0(GND), .Q1(GND), .Q2(GND) );

endmodule // dcntx4b

`endif

`ifdef dctlcar1
`else
`define dctlcar1
module dctlcar1( CLK , CLR, D, LOAD, Q, ACO1 );
output ACO1;
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [3:0] D;
input LOAD;
 input [3:0] Q;
wire N_1;
supply0 GND;
supply1 VCC;
wire N_2;
wire N_3;
wire N_4;
wire N_5;

dffp QL6 ( .CLK(CLK), .D(N_2), .PRE(CLR), .Q(ACO1) );
and4i3 QL5 ( .A(N_1), .B(LOAD), .C(Q[2]), .D(N_3), .Q(N_4) );
and4i3 QL4 ( .A(LOAD), .B(D[0]), .C(D[1]), .D(D[2]), .Q(N_5) );
dnflbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(VCC), .ENT(VCC), .LOAD(LOAD),
           .Q(N_3), .Q0(N_1), .Q1(GND), .Q2(GND) );
dnflbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(VCC), .ENT(VCC), .LOAD(LOAD),
           .Q(N_1), .Q0(GND), .Q1(GND), .Q2(GND) );
mux4x6 QL1 ( .A(GND), .B(Q[3]), .C(D[3]), .D(GND), .Q(N_2), .S0(N_4), .S1(N_5) );

endmodule // dctlcar1

`endif

`ifdef dcntl4c
`else
`define dcntl4c
module dcntl4c( CLK , CLR, D, ENP, ENT, LOAD, Q );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [3:0] D;
input ENP, ENT, LOAD;
 output [3:0] Q;
supply0 GND;

dnflbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
dnflbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(GND) );
dnflbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[1]), .Q0(Q[0]), .Q1(GND), .Q2(GND) );
dnflbit QL1 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[0]), .Q0(GND), .Q1(GND), .Q2(GND) );

endmodule // dcntl4c

`endif

`ifdef dctlcar3
`else
`define dctlcar3
module dctlcar3( CLK , CLR, D, LOAD, ACO1, ACO2, ACO3 );
output ACO1, ACO2, ACO3;
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [1:0] D;
input LOAD;
supply0 GND;
supply1 VCC;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;
wire N_9;
wire N_10;
wire N_11;

dffp QL14 ( .CLK(CLK), .D(N_3), .PRE(CLR), .Q(ACO3) );
dffp QL13 ( .CLK(CLK), .D(N_2), .PRE(CLR), .Q(ACO2) );
dffp QL12 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO1) );
and3i2 QL11 ( .A(LOAD), .B(D[0]), .C(D[1]), .Q(N_9) );
and3i2 QL10 ( .A(N_4), .B(N_5), .C(LOAD), .Q(N_6) );
and3i2 QL9 ( .A(LOAD), .B(D[0]), .C(D[1]), .Q(N_10) );
and3i2 QL8 ( .A(N_4), .B(N_5), .C(LOAD), .Q(N_7) );
and3i2 QL7 ( .A(LOAD), .B(D[0]), .C(D[1]), .Q(N_11) );
and3i2 QL6 ( .A(N_4), .B(N_5), .C(LOAD), .Q(N_8) );
dnflbit QL5 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(VCC), .ENT(VCC), .LOAD(LOAD),
           .Q(N_5), .Q0(N_4), .Q1(GND), .Q2(GND) );
dnflbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(VCC), .ENT(VCC), .LOAD(LOAD),
           .Q(N_4), .Q0(GND), .Q1(GND), .Q2(GND) );
mux4x0 QL3 ( .A(GND), .B(VCC), .C(VCC), .D(GND), .Q(N_1), .S0(N_6), .S1(N_9) );
mux4x0 QL2 ( .A(GND), .B(VCC), .C(VCC), .D(GND), .Q(N_2), .S0(N_7), .S1(N_10) );
mux4x0 QL1 ( .A(GND), .B(VCC), .C(VCC), .D(GND), .Q(N_3), .S0(N_8), .S1(N_11) );

endmodule // dctlcar3

`endif

`ifdef dctlcar2
`else
`define dctlcar2
module dctlcar2( CLK , CLR, D, LOAD, ACO1, ACO2 );
output ACO1, ACO2;
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [1:0] D;
input LOAD;
supply0 GND;
supply1 VCC;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
wire N_5;
wire N_6;
wire N_7;
wire N_8;

dffp QL10 ( .CLK(CLK), .D(N_2), .PRE(CLR), .Q(ACO2) );
dffp QL9 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO1) );
and3i2 QL8 ( .A(LOAD), .B(D[0]), .C(D[1]), .Q(N_7) );
and3i2 QL7 ( .A(N_3), .B(N_4), .C(LOAD), .Q(N_5) );
and3i2 QL6 ( .A(N_3), .B(N_4), .C(LOAD), .Q(N_6) );
and3i2 QL5 ( .A(LOAD), .B(D[0]), .C(D[1]), .Q(N_8) );
dnflbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(VCC), .ENT(VCC), .LOAD(LOAD),
           .Q(N_4), .Q0(N_3), .Q1(GND), .Q2(GND) );
dnflbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(VCC), .ENT(VCC), .LOAD(LOAD),
           .Q(N_3), .Q0(GND), .Q1(GND), .Q2(GND) );
mux4x0 QL2 ( .A(GND), .B(VCC), .C(VCC), .D(GND), .Q(N_1), .S0(N_5), .S1(N_7) );
mux4x0 QL1 ( .A(GND), .B(VCC), .C(VCC), .D(GND), .Q(N_2), .S0(N_6), .S1(N_8) );

endmodule // dctlcar2

`endif

`ifdef dcntl4b
`else
`define dcntl4b
module dcntl4b( CLK , CLR, D, ENP, ENT, LOAD, Q, RCO );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [3:0] D;
input ENP, ENT, LOAD;
 output [3:0] Q;
output RCO;
supply0 GND;

and5i4 QL5 ( .A(ENT), .B(Q[0]), .C(Q[1]), .D(Q[2]), .E(Q[3]), .Q(RCO) );
dnflbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
dnflbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(GND) );
dnflbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[1]), .Q0(Q[0]), .Q1(GND), .Q2(GND) );
dnflbit QL1 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(ENP), .ENT(ENT), .LOAD(LOAD),
           .Q(Q[0]), .Q0(GND), .Q1(GND), .Q2(GND) );

endmodule // dcntl4b

`endif

`ifdef dcntl4a
`else
`define dcntl4a
module dcntl4a( CLK , CLR, D, LOAD, Q, RCO );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
 input [3:0] D;
input LOAD;
 output [3:0] Q;
output RCO;
supply0 GND;
supply1 VCC;

and2i2 QL5 ( .A(Q[2]), .B(Q[3]), .Q(RCO) );
dnflbit QL4 ( .CLK(CLK), .CLR(CLR), .D(D[3]), .ENP(VCC), .ENT(VCC), .LOAD(LOAD),
           .Q(Q[3]), .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
dnflbit QL3 ( .CLK(CLK), .CLR(CLR), .D(D[2]), .ENP(VCC), .ENT(VCC), .LOAD(LOAD),
           .Q(Q[2]), .Q0(Q[0]), .Q1(Q[1]), .Q2(GND) );
dnflbit QL2 ( .CLK(CLK), .CLR(CLR), .D(D[1]), .ENP(VCC), .ENT(VCC), .LOAD(LOAD),
           .Q(Q[1]), .Q0(Q[0]), .Q1(GND), .Q2(GND) );
dnflbit QL1 ( .CLK(CLK), .CLR(CLR), .D(D[0]), .ENP(VCC), .ENT(VCC), .LOAD(LOAD),
           .Q(Q[0]), .Q0(GND), .Q1(GND), .Q2(GND) );

endmodule // dcntl4a

`endif

`ifdef dctecar1
`else
`define dctecar1
module dctecar1( CLK , CLR, ENG, Q, ACO1 );
output ACO1;
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input ENG;
 input [3:0] Q;
supply0 GND;
supply1 VCC;
wire N_1;
wire N_2;
wire N_3;
wire N_4;

dffp QL5 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO1) );
mux4x2 QL4 ( .A(GND), .B(N_3), .C(GND), .D(N_3), .Q(N_1), .S0(N_2), .S1(ENG) );
and3i3 QL3 ( .A(N_4), .B(Q[2]), .C(Q[3]), .Q(N_2) );
dnfebit QL2 ( .CLK(CLK), .CLR(CLR), .ENG(VCC), .ENP(ENG), .ENT(VCC), .Q(N_4),
           .Q0(N_3), .Q1(GND), .Q2(GND) );
dnfebit QL1 ( .CLK(CLK), .CLR(CLR), .ENG(VCC), .ENP(ENG), .ENT(VCC), .Q(N_3),
           .Q0(GND), .Q1(GND), .Q2(GND) );

endmodule // dctecar1

`endif

`ifdef dcnte4c
`else
`define dcnte4c
module dcnte4c( CLK , CLR, ENG, ENP, ENT, Q );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input ENG, ENP, ENT;
 output [3:0] Q;
supply0 GND;

dnfebit QL4 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(ENP), .ENT(ENT), .Q(Q[3]),
           .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
dnfebit QL3 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(ENP), .ENT(ENT), .Q(Q[2]),
           .Q0(Q[0]), .Q1(Q[1]), .Q2(GND) );
dnfebit QL2 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(ENP), .ENT(ENT), .Q(Q[1]),
           .Q0(Q[0]), .Q1(GND), .Q2(GND) );
dnfebit QL1 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(ENP), .ENT(ENT), .Q(Q[0]),
           .Q0(GND), .Q1(GND), .Q2(GND) );

endmodule // dcnte4c

`endif

`ifdef dcnte4b
`else
`define dcnte4b
module dcnte4b( CLK , CLR, ENG, ENP, ENT, Q, RCO );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input ENG, ENP, ENT;
 output [3:0] Q;
output RCO;
supply0 GND;

and5i4 QL5 ( .A(ENT), .B(Q[0]), .C(Q[1]), .D(Q[2]), .E(Q[3]), .Q(RCO) );
dnfebit QL4 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(ENP), .ENT(ENT), .Q(Q[3]),
           .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
dnfebit QL3 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(ENP), .ENT(ENT), .Q(Q[2]),
           .Q0(Q[0]), .Q1(Q[1]), .Q2(GND) );
dnfebit QL2 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(ENP), .ENT(ENT), .Q(Q[1]),
           .Q0(Q[0]), .Q1(GND), .Q2(GND) );
dnfebit QL1 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(ENP), .ENT(ENT), .Q(Q[0]),
           .Q0(GND), .Q1(GND), .Q2(GND) );

endmodule // dcnte4b

`endif

`ifdef dcnte4a
`else
`define dcnte4a
module dcnte4a( CLK , CLR, ENG, Q, RCO );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input ENG;
 output [3:0] Q;
output RCO;
supply1 VCC;
supply0 GND;

dnfebit QL1 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(VCC), .ENT(VCC), .Q(Q[0]),
           .Q0(GND), .Q1(GND), .Q2(GND) );
dnfebit QL2 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(VCC), .ENT(VCC), .Q(Q[1]),
           .Q0(Q[0]), .Q1(GND), .Q2(GND) );
dnfebit QL3 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(VCC), .ENT(VCC), .Q(Q[2]),
           .Q0(Q[0]), .Q1(Q[1]), .Q2(GND) );
dnfebit QL4 ( .CLK(CLK), .CLR(CLR), .ENG(ENG), .ENP(VCC), .ENT(VCC), .Q(Q[3]),
           .Q0(Q[0]), .Q1(Q[1]), .Q2(Q[2]) );
and2i2 QL5 ( .A(Q[2]), .B(Q[3]), .Q(RCO) );

endmodule // dcnte4a

`endif

`ifdef dnfecar3
`else
`define dnfecar3
module dnfecar3( CLK , CLR, ENG, ACO1, ACO2, ACO3 );
output ACO1, ACO2, ACO3;
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input ENG;
wire N_1;
wire N_2;
wire N_3;
wire N_4;
supply1 VCC;
supply0 GND;
wire N_5;

mux4x1 QL1 ( .A(N_4), .B(GND), .C(N_4), .D(GND), .Q(N_5), .S0(N_1), .S1(ENG) );
mux4x1 QL2 ( .A(N_4), .B(GND), .C(N_4), .D(GND), .Q(N_3), .S0(N_1), .S1(ENG) );
mux4x1 QL3 ( .A(N_4), .B(GND), .C(N_4), .D(GND), .Q(N_2), .S0(N_1), .S1(ENG) );
dnfebit QL4 ( .CLK(CLK), .CLR(CLR), .ENG(VCC), .ENP(ENG), .ENT(VCC), .Q(N_4),
           .Q0(GND), .Q1(GND), .Q2(GND) );
dnfebit QL5 ( .CLK(CLK), .CLR(CLR), .ENG(VCC), .ENP(ENG), .ENT(VCC), .Q(N_1),
           .Q0(N_4), .Q1(GND), .Q2(GND) );
dffp QL6 ( .CLK(CLK), .D(N_3), .PRE(CLR), .Q(ACO2) );
dffp QL7 ( .CLK(CLK), .D(N_2), .PRE(CLR), .Q(ACO3) );
dffp QL8 ( .CLK(CLK), .D(N_5), .PRE(CLR), .Q(ACO1) );

endmodule // dnfecar3

`endif

`ifdef dnfecar2
`else
`define dnfecar2
module dnfecar2( CLK , CLR, ENG, ACO1, ACO2 );
output ACO1, ACO2;
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input ENG;
supply1 VCC;
supply0 GND;
wire N_1;
wire N_2;
wire N_3;
wire N_4;

dffp QL6 ( .CLK(CLK), .D(N_2), .PRE(CLR), .Q(ACO2) );
dffp QL5 ( .CLK(CLK), .D(N_1), .PRE(CLR), .Q(ACO1) );
mux4x1 QL4 ( .A(N_3), .B(GND), .C(N_3), .D(GND), .Q(N_2), .S0(N_4), .S1(ENG) );
mux4x1 QL3 ( .A(N_3), .B(GND), .C(N_3), .D(GND), .Q(N_1), .S0(N_4), .S1(ENG) );
dnfebit QL2 ( .CLK(CLK), .CLR(CLR), .ENG(VCC), .ENP(ENG), .ENT(VCC), .Q(N_4),
           .Q0(N_3), .Q1(GND), .Q2(GND) );
dnfebit QL1 ( .CLK(CLK), .CLR(CLR), .ENG(VCC), .ENP(ENG), .ENT(VCC), .Q(N_3),
           .Q0(GND), .Q1(GND), .Q2(GND) );

endmodule // dnfecar2

`endif

`ifdef csamuxa
`else
`define csamuxa
module csamuxa( A , S00, S01, S1, Q );
input A;
output Q;
input S00, S01, S1;

mux4xa QL1 ( .A(S00), .B(S00), .C(S01), .D(S01), .Q(Q), .S0(A), .S1(S1) );

endmodule // csamuxa

`endif

`ifdef csamuxb
`else
`define csamuxb
module csamuxb( A , B, S00, S01, S1, Q );
input A, B;
output Q;
input S00, S01, S1;
wire N_1;

and2i0 QL1 ( .A(S1), .B(S01), .Q(N_1) );
mux4x0 QL2 ( .A(A), .B(B), .C(B), .D(B), .Q(Q), .S0(N_1), .S1(S00) );

endmodule // csamuxb

`endif

`ifdef csamuxc
`else
`define csamuxc
module csamuxc( A , B, S00, S01, S1, Q );
input A, B;
output Q;
input S00, S01, S1;
wire N_1;

and2i1 QL1 ( .A(S1), .B(S01), .Q(N_1) );
mux4xe QL2 ( .A(A), .B(B), .C(B), .D(B), .Q(Q), .S0(N_1), .S1(S00) );

endmodule // csamuxc

`endif

`ifdef csamuxd
`else
`define csamuxd
module csamuxd( A , S00, S01, S1, Q );
input A;
output Q;
input S00, S01, S1;

mux4x6 QL1 ( .A(S00), .B(S00), .C(S01), .D(S01), .Q(Q), .S0(A), .S1(S1) );

endmodule // csamuxd

`endif

`ifdef muxb2dx2
`else
`define muxb2dx2
module muxb2dx2( A , B, C, D, S, Q, R, T );
input A, B, C, D;
output Q, R;
input S;
output T;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
supply1 VCC;

frag_m I_2 ( .B1(A), .B2(GND), .C1(VCC), .C2(B), .D1(C), .D2(GND), .E1(VCC), .E2(D),
          .NS(T), .NZ(R), .OS(N_1), .OZ(Q) );
frag_f I_1 ( .F1(S), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(T) );
frag_a QL1 ( .A1(GND), .A2(VCC), .A3(GND), .A4(VCC), .A5(GND), .A6(VCC), .AZ(N_1) );

endmodule // muxb2dx2

`endif

`ifdef muxc2dx2
`else
`define muxc2dx2
module muxc2dx2( A , B, C, D, S, Q, R, T );
input A, B, C, D;
output Q, R;
input S;
output T;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
supply1 VCC;

frag_m I_2 ( .B1(VCC), .B2(B), .C1(A), .C2(GND), .D1(VCC), .D2(D), .E1(C), .E2(GND),
          .NS(T), .NZ(R), .OS(N_1), .OZ(Q) );
frag_f I_1 ( .F1(S), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(T) );
frag_a QL1 ( .A1(GND), .A2(VCC), .A3(GND), .A4(VCC), .A5(GND), .A6(VCC), .AZ(N_1) );

endmodule // muxc2dx2

`endif

`ifdef xor2p
`else
`define xor2p
module xor2p( A , B, Q );
input A, B;
output Q;
supply1 VCC;
supply0 GND;

mux4x0 QL1 ( .A(GND), .B(VCC), .C(VCC), .D(GND), .Q(Q), .S0(B), .S1(A) );

endmodule // xor2p

`endif

`ifdef csblow
`else
`define csblow
module csblow( A0 , A1, B0, B1, A1T, C0_n, C1 );
input A0, A1;
output A1T;
input B0, B1;
output C0_n, C1;
parameter ql_gate = `LOGIC;
supply0 GND;
supply1 VCC;

frag_m I_2 ( .B1(VCC), .B2(B1), .C1(VCC), .C2(GND), .D1(GND), .D2(VCC), .E1(VCC),
          .E2(B1), .NS(A1T), .OS(C0_n), .OZ(C1) );
frag_f I_1 ( .F1(A1), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(A1T) );
frag_a QL1 ( .A1(VCC), .A2(A0), .A3(B0), .A4(GND), .A5(VCC), .A6(GND), .AZ(C0_n) );

endmodule // csblow

`endif

`ifdef csbbitb
`else
`define csbbitb
module csbbitb( A , B, C0, C1, S0 );
input A, B;
output C0, C1, S0;
parameter ql_gate = `LOGIC;
supply0 GND;
supply1 VCC;

frag_m I_2 ( .B1(VCC), .B2(GND), .C1(GND), .C2(VCC), .D1(GND), .D2(VCC), .E1(GND),
          .E2(VCC), .NS(C1), .OS(C0), .OZ(S0) );
frag_f I_1 ( .F1(VCC), .F2(GND), .F3(VCC), .F4(GND), .F5(B), .F6(A), .FZ(C1) );
frag_a QL1 ( .A1(A), .A2(GND), .A3(VCC), .A4(B), .A5(VCC), .A6(GND), .AZ(C0) );

endmodule // csbbitb

`endif

`ifdef csbbita
`else
`define csbbita
module csbbita( A , B, C0, C1, S0 );
input A, B;
output C0, C1, S0;

and2i2 QL1 ( .A(C0), .B(C1), .Q(S0) );
nor2i1 QL2 ( .A(A), .B(B), .Q(C1) );
and2i1 QL3 ( .A(A), .B(B), .Q(C0) );

endmodule // csbbita

`endif

`ifdef mux2dxy
`else
`define mux2dxy
module mux2dxy( A , B, C, D, S, Q, R );
input A, B, C, D;
output Q, R;
input S;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply0 GND;
supply1 VCC;

frag_m I_2 ( .B1(A), .B2(GND), .C1(VCC), .C2(B), .D1(VCC), .D2(C), .E1(D), .E2(GND),
          .NS(N_1), .NZ(R), .OS(N_2), .OZ(Q) );
frag_f I_1 ( .F1(S), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_a QL1 ( .A1(GND), .A2(VCC), .A3(GND), .A4(VCC), .A5(GND), .A6(VCC), .AZ(N_2) );

endmodule // mux2dxy

`endif

`ifdef xnor2p
`else
`define xnor2p
module xnor2p( A , B, Q );
input A, B;
output Q;
supply1 VCC;
supply0 GND;

mux4x0 QL1 ( .A(VCC), .B(GND), .C(GND), .D(VCC), .Q(Q), .S0(B), .S1(A) );

endmodule // xnor2p

`endif

`ifdef muxb2dx0
`else
`define muxb2dx0
module muxb2dx0( A , B, C, D, S, Q, R, T );
input A, B, C, D;
output Q, R;
input S;
output T;
parameter ql_gate = `LOGIC;
wire N_1;
supply0 GND;
supply1 VCC;

frag_m I_2 ( .B1(A), .B2(GND), .C1(B), .C2(GND), .D1(C), .D2(GND), .E1(D), .E2(GND),
          .NS(T), .NZ(R), .OS(N_1), .OZ(Q) );
frag_f I_1 ( .F1(S), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(T) );
frag_a QL1 ( .A1(GND), .A2(VCC), .A3(GND), .A4(VCC), .A5(GND), .A6(VCC), .AZ(N_1) );

endmodule // muxb2dx0

`endif

`ifdef mux2dxx
`else
`define mux2dxx
module mux2dxx( A , B, C, D, S, Q, R );
input A, B, C, D;
output Q, R;
input S;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply0 GND;
supply1 VCC;

frag_m I_2 ( .B1(A), .B2(GND), .C1(VCC), .C2(B), .D1(C), .D2(GND), .E1(D), .E2(GND),
          .NS(N_1), .NZ(R), .OS(N_2), .OZ(Q) );
frag_f I_1 ( .F1(S), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_1) );
frag_a QL1 ( .A1(GND), .A2(VCC), .A3(GND), .A4(VCC), .A5(GND), .A6(VCC), .AZ(N_2) );

endmodule // mux2dxx

`endif

`ifdef muxi2dx2
`else
`define muxi2dx2
module muxi2dx2( A , B, C, D, S, Q, R );
input A, B, C, D;
output Q, R;
input S;

mux2dx1 QL1 ( .A(B), .B(A), .C(D), .D(C), .Q(Q), .R(R), .S(S) );

endmodule // muxi2dx2

`endif

`ifdef mbitc
`else
`define mbitc
module mbitc( A , B0, B1, CI, CO, S );
input A, B0, B1, CI;
output CO, S;
wire N_1;
wire N_2;

maj3i0 QL4 ( .A(A), .B(N_2), .C(CI), .Q(CO) );
and2i0 QL3 ( .A(B0), .B(B1), .Q(N_2) );
and2i0 QL2 ( .A(B0), .B(B1), .Q(N_1) );
xor3i0 QL1 ( .A(A), .B(N_1), .C(CI), .Q(S) );

endmodule // mbitc

`endif

`ifdef mbitb
`else
`define mbitb
module mbitb( A0 , A1, B, CI, CO, S );
input A0, A1, B, CI;
output CO, S;
wire N_1;
wire N_2;

maj3i0 QL1 ( .A(N_1), .B(B), .C(CI), .Q(CO) );
and2i0 QL2 ( .A(A0), .B(A1), .Q(N_1) );
and2i0 QL3 ( .A(A0), .B(A1), .Q(N_2) );
xor3i0 QL4 ( .A(N_2), .B(B), .C(CI), .Q(S) );

endmodule // mbitb

`endif

`ifdef mbita
`else
`define mbita
module mbita( A0 , A1, B0, B1, CI, CO, S );
input A0, A1, B0, B1, CI;
output CO, S;
wire N_1;
wire N_2;
wire N_3;
wire N_4;

xor3i0 QL1 ( .A(N_2), .B(N_4), .C(CI), .Q(S) );
and2i0 QL2 ( .A(A0), .B(A1), .Q(N_1) );
and2i0 QL3 ( .A(B0), .B(B1), .Q(N_4) );
and2i0 QL4 ( .A(A0), .B(A1), .Q(N_2) );
and2i0 QL5 ( .A(B0), .B(B1), .Q(N_3) );
maj3i0 QL6 ( .A(N_1), .B(N_3), .C(CI), .Q(CO) );

endmodule // mbita

`endif

`ifdef eqcombit
`else
`define eqcombit
module eqcombit( A1 , A2, B1, B2, EQ1, EQ2 );
input A1, A2, B1, B2;
output EQ1, EQ2;
parameter syn_macro = 1, ql_pack = 1;
parameter ql_gate = `LOGIC;
supply0 GND;
supply1 VCC;
wire N_1;
wire N_2;

frag_m I_2 ( .B1(B1), .B2(A1), .C1(B1), .C2(A1), .D1(VCC), .D2(A2), .E1(A2),
          .E2(GND), .NS(N_2), .NZ(EQ2), .OS(N_1), .OZ(EQ1) );
frag_f I_1 ( .F1(B2), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(N_2) );
frag_a QL1 ( .A1(A1), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(B1), .AZ(N_1) );

endmodule // eqcombit

`endif

`ifdef csalow
`else
`define csalow
module csalow( A0 , A1, B0, B1, A1T, C0, C1 );
input A0, A1;
output A1T;
input B0, B1;
output C0, C1;
parameter ql_gate = `LOGIC;
supply0 GND;
supply1 VCC;

frag_m I_2 ( .B1(GND), .B2(VCC), .C1(B1), .C2(GND), .D1(B1), .D2(GND), .E1(VCC),
          .E2(GND), .NS(A1T), .OS(C0), .OZ(C1) );
frag_f I_1 ( .F1(A1), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GND), .FZ(A1T) );
frag_a QL1 ( .A1(A0), .A2(GND), .A3(B0), .A4(GND), .A5(VCC), .A6(GND), .AZ(C0) );

endmodule // csalow

`endif

`ifdef csabita
`else
`define csabita
module csabita( A , B, C0, C1, S0 );
input A, B;
output C0, C1, S0;

and2i0 QL1 ( .A(A), .B(B), .Q(C0) );
nor2i0 QL2 ( .A(A), .B(B), .Q(C1) );
and2i2 QL3 ( .A(C0), .B(C1), .Q(S0) );

endmodule // csabita

`endif

`ifdef csabitb
`else
`define csabitb
module csabitb( A , B, C0, C1, S0 );
input A, B;
output C0, C1, S0;
parameter ql_gate = `LOGIC;
supply0 GND;
supply1 VCC;

frag_m I_2 ( .B1(VCC), .B2(GND), .C1(GND), .C2(VCC), .D1(GND), .D2(VCC), .E1(GND),
          .E2(VCC), .NS(C1), .OS(C0), .OZ(S0) );
frag_f I_1 ( .F1(VCC), .F2(GND), .F3(VCC), .F4(B), .F5(VCC), .F6(A), .FZ(C1) );
frag_a QL1 ( .A1(A), .A2(GND), .A3(B), .A4(GND), .A5(VCC), .A6(GND), .AZ(C0) );

endmodule // csabitb

`endif

`ifdef upflbit
`else
`define upflbit
module upflbit( CLK , CLR, D, ENP, ENT, LOAD, Q0, Q1, Q2, Q );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input D, ENP, ENT, LOAD;
output Q;
input Q0, Q1, Q2;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(GND), .QZ(Q) );
frag_m I_2 ( .B1(D), .B2(GND), .C1(D), .C2(GND), .D1(Q), .D2(GND), .E1(VCC), .E2(Q),
          .NS(N_2), .OS(N_3), .OZ(N_1) );
frag_f I_1 ( .F1(Q0), .F2(ENP), .F3(Q1), .F4(ENT), .F5(Q2), .F6(GND), .FZ(N_2) );
frag_a QL1 ( .A1(LOAD), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_3) );

endmodule // upflbit

`endif

`ifdef upfxbit
`else
`define upfxbit
module upfxbit( CLK , CLR, D, ENG, ENP, ENT, LOAD, Q0, Q1, Q2, Q );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input D, ENG, ENP, ENT, LOAD;
output Q;
input Q0, Q1, Q2;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(GND), .QZ(Q) );
frag_m I_2 ( .B1(Q), .B2(GND), .C1(VCC), .C2(Q), .D1(D), .D2(GND), .E1(D), .E2(GND),
          .NS(N_2), .OS(N_3), .OZ(N_1) );
frag_f I_1 ( .F1(Q0), .F2(ENP), .F3(Q1), .F4(ENT), .F5(Q2), .F6(ENG), .FZ(N_2) );
frag_a QL1 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(LOAD), .AZ(N_3) );

endmodule // upfxbit

`endif

`ifdef borrow0
`else
`define borrow0
module borrow0( A , B, Bin, Bout );
input A, B, Bin;
output Bout;
parameter ql_gate = `LOGIC;
supply1 vcc;
supply0 GNd;

lcell2 I_3 ( .A1(vcc), .A2(Bin), .A3(vcc), .A4(GNd), .A5(vcc), .A6(GNd), .B1(GNd),
          .B2(GNd), .C1(vcc), .C2(B), .D1(A), .D2(GNd), .E1(vcc), .E2(GNd),
          .F1(vcc), .F2(B), .F3(vcc), .F4(GNd), .F5(vcc), .F6(GNd), .MP(GNd),
          .MS(A), .NP(vcc), .NS(GNd), .OP(vcc), .OS(GNd), .OZ(Bout), .QC(GNd),
          .QR(GNd), .QS(GNd) );

endmodule // borrow0

`endif

`ifdef dif0
`else
`define dif0
module dif0( A , B, Bin, d0 );
input A, B, Bin;
output d0;
parameter ql_gate = `LOGIC;
supply1 vcc;
supply0 gnd;

lcell2 I_3 ( .A1(vcc), .A2(Bin), .A3(vcc), .A4(gnd), .A5(vcc), .A6(gnd), .B1(vcc),
          .B2(A), .C1(A), .C2(gnd), .D1(B), .D2(gnd), .E1(vcc), .E2(B), .F1(gnd),
          .F2(gnd), .F3(gnd), .F4(gnd), .F5(gnd), .F6(gnd), .MP(gnd), .MS(B),
          .NP(gnd), .NS(A), .OP(vcc), .OS(gnd), .OZ(d0), .QC(gnd), .QR(gnd),
          .QS(gnd) );

endmodule // dif0

`endif

`ifdef sum2_gen
`else
`define sum2_gen
module sum2_gen( C_i , Cj_i0, Cj_i1, Ck_j0, Ck_j1, Sk_0, Sk_1, Sk_i );
input C_i, Cj_i0, Cj_i1, Ck_j0, Ck_j1, Sk_0, Sk_1;
output Sk_i;
parameter ql_gate = `LOGIC;
supply0 gnd;
supply1 vcc;

lcell2 I_3 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(Cj_i1), .A6(gnd),
          .B1(Sk_0), .B2(gnd), .C1(Sk_1), .C2(gnd), .D1(Sk_0), .D2(gnd),
          .E1(Sk_1), .E2(gnd), .F1(gnd), .F2(gnd), .F3(gnd), .F4(gnd), .F5(gnd),
          .F6(gnd), .MP(gnd), .MS(Ck_j0), .NP(gnd), .NS(Ck_j1), .OP(C_i),
          .OS(Cj_i0), .OZ(Sk_i), .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // sum2_gen

`endif

`ifdef cary_gen
`else
`define cary_gen
module cary_gen( C_i , Cj_i0, Cj_i1, Ck_j0, Ck_j1, Cm_k0, Cm_k1, Cm_i );
input C_i, Cj_i0, Cj_i1, Ck_j0, Ck_j1;
output Cm_i;
input Cm_k0, Cm_k1;
parameter ql_gate = `LOGIC;
supply0 gnd;
supply1 vcc;

lcell2 I_3 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(Cj_i1), .A6(gnd),
          .B1(Cm_k0), .B2(gnd), .C1(Cm_k1), .C2(gnd), .D1(Cm_k0), .D2(gnd),
          .E1(Cm_k1), .E2(gnd), .F1(gnd), .F2(gnd), .F3(gnd), .F4(gnd), .F5(gnd),
          .F6(gnd), .MP(gnd), .MS(Ck_j0), .NP(gnd), .NS(Ck_j1), .OP(C_i),
          .OS(Cj_i0), .OZ(Cm_i), .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // cary_gen

`endif

`ifdef sum_gen
`else
`define sum_gen
module sum_gen( C_i , Cj_i0, Cj_i1, Ck_j0, Ck_j1, Sk_01, Sk_i );
input C_i, Cj_i0, Cj_i1, Ck_j0, Ck_j1, Sk_01;
output Sk_i;
parameter ql_gate = `LOGIC;
supply0 gnd;
supply1 vcc;

lcell2 I_3 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(Cj_i1), .A6(gnd),
          .B1(Sk_01), .B2(gnd), .C1(vcc), .C2(Sk_01), .D1(Sk_01), .D2(gnd),
          .E1(vcc), .E2(Sk_01), .F1(gnd), .F2(gnd), .F3(gnd), .F4(gnd), .F5(gnd),
          .F6(gnd), .MP(gnd), .MS(Ck_j0), .NP(gnd), .NS(Ck_j1), .OP(C_i),
          .OS(Cj_i0), .OZ(Sk_i), .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // sum_gen

`endif

`ifdef dif_b0
`else
`define dif_b0
module dif_b0( Ax , Bx, Bo_Bi0, Bo_Bi1 );
input Ax;
output Bo_Bi0, Bo_Bi1;
input Bx;
parameter ql_gate = `LOGIC;
supply1 vcc;
supply0 gnd;

lcell2 I_3 ( .A1(gnd), .A2(gnd), .A3(gnd), .A4(gnd), .A5(gnd), .A6(gnd), .B1(vcc),
          .B2(Bx), .C1(vcc), .C2(gnd), .D1(vcc), .D2(Bx), .E1(Bx), .E2(gnd),
          .F1(Ax), .F2(gnd), .F3(vcc), .F4(Bx), .F5(vcc), .F6(gnd), .FZ(Bo_Bi0),
          .MP(gnd), .MS(Ax), .NP(gnd), .NS(Ax), .OP(gnd), .OS(gnd), .OZ(Bo_Bi1),
          .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // dif_b0

`endif

`ifdef dif_b
`else
`define dif_b
module dif_b( Ax , Bx, Bo_Bi0, Bo_Bi1, Sub_Dif );
input Ax;
output Bo_Bi0, Bo_Bi1;
input Bx;
output Sub_Dif;
parameter ql_gate = `LOGIC;
supply1 vcc;
supply0 gnd;

lcell2 I_3 ( .A1(gnd), .A2(gnd), .A3(gnd), .A4(gnd), .A5(gnd), .A6(gnd), .B1(vcc),
          .B2(Bx), .C1(vcc), .C2(gnd), .D1(vcc), .D2(Bx), .E1(Bx), .E2(gnd),
          .F1(Ax), .F2(gnd), .F3(vcc), .F4(Bx), .F5(vcc), .F6(gnd), .FZ(Bo_Bi0),
          .MP(gnd), .MS(Ax), .NP(gnd), .NS(Ax), .NZ(Sub_Dif), .OP(gnd), .OS(gnd),
          .OZ(Bo_Bi1), .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // dif_b

`endif

`ifdef b_out
`else
`define b_out
module b_out( By_x0 , Bz_y0, Bz_y1, Bo );
output Bo;
input By_x0, Bz_y0, Bz_y1;
parameter ql_gate = `LOGIC;
supply0 gnd;
supply1 vcc;

lcell2 I_3 ( .A1(gnd), .A2(gnd), .A3(gnd), .A4(gnd), .A5(gnd), .A6(gnd), .B1(vcc),
          .B2(Bz_y0), .C1(vcc), .C2(Bz_y1), .D1(gnd), .D2(gnd), .E1(gnd),
          .E2(gnd), .F1(gnd), .F2(gnd), .F3(gnd), .F4(gnd), .F5(gnd), .F6(gnd),
          .MP(gnd), .MS(By_x0), .NP(gnd), .NS(gnd), .OP(gnd), .OS(gnd), .OZ(Bo),
          .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // b_out

`endif

`ifdef bo_gen
`else
`define bo_gen
module bo_gen( C_i , Cj_i0, Cj_i1, Ck_j0, Ck_j1, Cm_k0, Cm_k1, Cm_i );
input C_i, Cj_i0, Cj_i1, Ck_j0, Ck_j1;
output Cm_i;
input Cm_k0, Cm_k1;
parameter ql_gate = `LOGIC;
supply0 gnd;
supply1 vcc;

lcell2 I_3 ( .A1(vcc), .A2(gnd), .A3(vcc), .A4(gnd), .A5(Cj_i1), .A6(gnd), .B1(vcc),
          .B2(Cm_k0), .C1(vcc), .C2(Cm_k1), .D1(vcc), .D2(Cm_k0), .E1(vcc),
          .E2(Cm_k1), .F1(gnd), .F2(gnd), .F3(gnd), .F4(gnd), .F5(gnd), .F6(gnd),
          .MP(gnd), .MS(Ck_j0), .NP(gnd), .NS(Ck_j1), .OP(C_i), .OS(Cj_i0),
          .OZ(Cm_i), .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // bo_gen

`endif

`ifdef sum_c0
`else
`define sum_c0
module sum_c0( Ax , Bx, Co_Ci0, Co_Ci1 );
input Ax, Bx;
output Co_Ci0, Co_Ci1;
parameter ql_gate = `LOGIC;
supply1 vcc;
supply0 gnd;

lcell2 I_3 ( .A1(gnd), .A2(gnd), .A3(gnd), .A4(gnd), .A5(gnd), .A6(gnd), .B1(Bx),
          .B2(gnd), .C1(vcc), .C2(gnd), .D1(Bx), .D2(gnd), .E1(vcc), .E2(Bx),
          .F1(Ax), .F2(gnd), .F3(Bx), .F4(gnd), .F5(vcc), .F6(gnd), .FZ(Co_Ci0),
          .MP(gnd), .MS(Ax), .NP(gnd), .NS(Ax), .OP(gnd), .OS(gnd), .OZ(Co_Ci1),
          .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // sum_c0

`endif

`ifdef sum_c
`else
`define sum_c
module sum_c( Ax , Bx, Co_Ci0, Co_Ci1, Sub_Sum );
input Ax, Bx;
output Co_Ci0, Co_Ci1, Sub_Sum;
parameter ql_gate = `LOGIC;
supply1 vcc;
supply0 gnd;

lcell2 I_3 ( .A1(gnd), .A2(gnd), .A3(gnd), .A4(gnd), .A5(gnd), .A6(gnd), .B1(Bx),
          .B2(gnd), .C1(vcc), .C2(gnd), .D1(Bx), .D2(gnd), .E1(vcc), .E2(Bx),
          .F1(Ax), .F2(gnd), .F3(Bx), .F4(gnd), .F5(vcc), .F6(gnd), .FZ(Co_Ci0),
          .MP(gnd), .MS(Ax), .NP(gnd), .NS(Ax), .NZ(Sub_Sum), .OP(gnd), .OS(gnd),
          .OZ(Co_Ci1), .QC(gnd), .QR(gnd), .QS(gnd) );

endmodule // sum_c

`endif

`ifdef carry0
`else
`define carry0
module carry0( A , B, Cin, Cout );
input A, B, Cin;
output Cout;
parameter ql_gate = `LOGIC;
supply1 vcc;
supply0 GNd;

lcell2 I_3 ( .A1(GNd), .A2(GNd), .A3(GNd), .A4(GNd), .A5(GNd), .A6(GNd), .B1(GNd),
          .B2(GNd), .C1(B), .C2(GNd), .D1(A), .D2(GNd), .E1(vcc), .E2(GNd),
          .F1(GNd), .F2(GNd), .F3(GNd), .F4(GNd), .F5(GNd), .F6(GNd), .MP(GNd),
          .MS(A), .NP(GNd), .NS(B), .OP(GNd), .OS(Cin), .OZ(Cout), .QC(GNd),
          .QR(GNd), .QS(GNd) );

endmodule // carry0

`endif

`ifdef sum0
`else
`define sum0
module sum0( A , B, Cin, s0 );
input A, B, Cin;
output s0;
parameter ql_gate = `LOGIC;
supply1 vcc;
supply0 gnd;

lcell2 I_3 ( .A1(gnd), .A2(gnd), .A3(gnd), .A4(gnd), .A5(gnd), .A6(gnd), .B1(A),
          .B2(gnd), .C1(vcc), .C2(A), .D1(vcc), .D2(B), .E1(B), .E2(gnd),
          .F1(gnd), .F2(gnd), .F3(gnd), .F4(gnd), .F5(gnd), .F6(gnd), .MP(gnd),
          .MS(B), .NP(gnd), .NS(A), .OP(gnd), .OS(Cin), .OZ(s0), .QC(gnd),
          .QR(gnd), .QS(gnd) );

endmodule // sum0

`endif

`ifdef ltch259
`else
`define ltch259
module ltch259( CLRNN , DATA, DECIN, GNN, Q );
input CLRNN, DATA, DECIN, GNN;
output Q;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;
wire N_1;
wire N_2;

frag_f I_2 ( .F1(DECIN), .F2(GND), .F3(VCC), .F4(GND), .F5(VCC), .F6(GNN), .FZ(N_1) );
frag_m I_1 ( .B1(GND), .B2(VCC), .C1(DECIN), .C2(GND), .D1(Q), .D2(GND), .E1(DATA),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(Q) );
frag_a QL1 ( .A1(CLRNN), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_2) );

endmodule // ltch259

`endif

`ifdef updnbitb
`else
`define updnbitb
module updnbitb( CLK , CLR, D0, D1, ENP, ENT, U0, U1, UP, Q );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input D0, D1, ENP, ENT;
output Q;
input U0, U1, UP;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(GND), .QZ(Q) );
frag_m I_2 ( .B1(Q), .B2(GND), .C1(VCC), .C2(Q), .D1(VCC), .D2(Q), .E1(VCC),
          .E2(GND), .NS(N_2), .OS(N_3), .OZ(N_1) );
frag_f I_1 ( .F1(ENP), .F2(ENT), .F3(UP), .F4(D0), .F5(VCC), .F6(D1), .FZ(N_2) );
frag_a QL1 ( .A1(ENP), .A2(ENT), .A3(U0), .A4(UP), .A5(U1), .A6(GND), .AZ(N_3) );

endmodule // updnbitb

`endif

`ifdef updncarb
`else
`define updncarb
module updncarb( ENT , Q0, Q1, Q2, UP, CO );
output CO;
input ENT, Q0, Q1, Q2, UP;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply0 GND;
supply1 VCC;

frag_m I_2 ( .B1(VCC), .B2(GND), .C1(ENT), .C2(GND), .D1(ENT), .D2(GND), .E1(VCC),
          .E2(GND), .NS(N_1), .OS(N_2), .OZ(CO) );
frag_f I_1 ( .F1(UP), .F2(Q0), .F3(VCC), .F4(Q1), .F5(VCC), .F6(Q2), .FZ(N_1) );
frag_a QL1 ( .A1(Q0), .A2(UP), .A3(Q1), .A4(GND), .A5(Q2), .A6(GND), .AZ(N_2) );

endmodule // updncarb

`endif

`ifdef updnbita
`else
`define updnbita
module updnbita( CLK , CLR, D0, D1, ENP, ENT, U0, U1, UP, Q );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input D0, D1, ENP, ENT;
output Q;
input U0, U1, UP;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(GND), .QZ(Q) );
frag_m I_2 ( .B1(Q), .B2(GND), .C1(VCC), .C2(Q), .D1(VCC), .D2(Q), .E1(VCC),
          .E2(GND), .NS(N_2), .OS(N_3), .OZ(N_1) );
frag_f I_1 ( .F1(ENT), .F2(ENP), .F3(UP), .F4(D0), .F5(VCC), .F6(D1), .FZ(N_2) );
frag_a QL1 ( .A1(ENT), .A2(ENP), .A3(U0), .A4(UP), .A5(U1), .A6(GND), .AZ(N_3) );

endmodule // updnbita

`endif

`ifdef updncara
`else
`define updncara
module updncara( ENT , Q0, Q1, Q2, UP, CO );
output CO;
input ENT, Q0, Q1, Q2, UP;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
supply0 GND;
supply1 VCC;

frag_m I_2 ( .B1(GND), .B2(VCC), .C1(ENT), .C2(GND), .D1(ENT), .D2(GND), .E1(GND),
          .E2(VCC), .NS(N_1), .OS(N_2), .OZ(CO) );
frag_f I_1 ( .F1(UP), .F2(Q0), .F3(VCC), .F4(Q1), .F5(VCC), .F6(Q2), .FZ(N_1) );
frag_a QL1 ( .A1(Q0), .A2(UP), .A3(Q1), .A4(GND), .A5(Q2), .A6(GND), .AZ(N_2) );

endmodule // updncara

`endif

`ifdef upfebit
`else
`define upfebit
module upfebit( CLK , CLR, ENG, ENP, ENT, Q0, Q1, Q2, Q );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input ENG, ENP, ENT;
output Q;
input Q0, Q1, Q2;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(GND), .QZ(Q) );
frag_m I_2 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(Q), .D2(GND), .E1(VCC),
          .E2(Q), .NS(N_2), .OS(N_3), .OZ(N_1) );
frag_f I_1 ( .F1(Q0), .F2(ENP), .F3(Q1), .F4(ENT), .F5(Q2), .F6(ENG), .FZ(N_2) );
frag_a QL1 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_3) );

endmodule // upfebit

`endif

`ifdef dnfxbit
`else
`define dnfxbit
module dnfxbit( CLK , CLR, D, ENG, ENP, ENT, LOAD, Q0, Q1, Q2, Q );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input D, ENG, ENP, ENT, LOAD;
output Q;
input Q0, Q1, Q2;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(GND), .QZ(Q) );
frag_m I_2 ( .B1(Q), .B2(GND), .C1(VCC), .C2(Q), .D1(D), .D2(GND), .E1(D), .E2(GND),
          .NS(N_2), .OS(N_3), .OZ(N_1) );
frag_f I_1 ( .F1(ENP), .F2(Q0), .F3(ENT), .F4(Q1), .F5(ENG), .F6(Q2), .FZ(N_2) );
frag_a QL1 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(LOAD), .A6(GND), .AZ(N_3) );

endmodule // dnfxbit

`endif

`ifdef dnflbit
`else
`define dnflbit
module dnflbit( CLK , CLR, D, ENP, ENT, LOAD, Q0, Q1, Q2, Q );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input D, ENP, ENT, LOAD;
output Q;
input Q0, Q1, Q2;
parameter ql_gate = `LOGIC;
supply1 VCC;
supply0 GND;
wire N_1;
wire N_2;
wire N_3;

frag_a QL1 ( .A1(VCC), .A2(LOAD), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_1) );
frag_f I_1 ( .F1(ENT), .F2(Q0), .F3(ENP), .F4(Q1), .F5(VCC), .F6(Q2), .FZ(N_2) );
frag_m I_2 ( .B1(D), .B2(GND), .C1(D), .C2(GND), .D1(Q), .D2(GND), .E1(VCC), .E2(Q),
          .NS(N_2), .OS(N_1), .OZ(N_3) );
frag_q I_3 ( .QC(CLK), .QD(N_3), .QR(CLR), .QS(GND), .QZ(Q) );

endmodule // dnflbit

`endif

`ifdef dnfebit
`else
`define dnfebit
module dnfebit( CLK , CLR, ENG, ENP, ENT, Q0, Q1, Q2, Q );
input CLK /* synthesis syn_isclock =1 */;
input CLR /* synthesis syn_isclock =1 */;
input ENG, ENP, ENT;
output Q;
input Q0, Q1, Q2;
parameter ql_gate = `LOGIC;
wire N_1;
wire N_2;
wire N_3;
supply0 GND;
supply1 VCC;

frag_q I_3 ( .QC(CLK), .QD(N_1), .QR(CLR), .QS(GND), .QZ(Q) );
frag_m I_2 ( .B1(VCC), .B2(GND), .C1(VCC), .C2(GND), .D1(Q), .D2(GND), .E1(VCC),
          .E2(Q), .NS(N_2), .OS(N_3), .OZ(N_1) );
frag_f I_1 ( .F1(ENP), .F2(Q0), .F3(ENT), .F4(Q1), .F5(ENG), .F6(Q2), .FZ(N_2) );
frag_a QL1 ( .A1(VCC), .A2(GND), .A3(VCC), .A4(GND), .A5(VCC), .A6(GND), .AZ(N_3) );

endmodule // dnfebit

`endif
