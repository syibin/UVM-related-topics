//------------------------------------------------------------
//   Copyright 2018 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//   
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//   
//       http://www.apache.org/licenses/LICENSE-2.0
//   
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------


const string s_alu_config_id = "alu_config";

class alu_agent_config extends uvm_object;
  `uvm_object_utils( alu_agent_config );

// Configuration Parameters
  virtual alu_monitor_bfm mon_bfm;
  virtual alu_driver_bfm  drv_bfm;
  int lock_num;
  string alu_seqr_name;


// Methods
  function new( string name = "alu_agent_config" );
    super.new( name );
  endfunction

endclass

