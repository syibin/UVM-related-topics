`define APB_FSM_IDLE 0
`define APB_FSM_SETUP 1
`define APB_FSM_ACCESS 2
`define APB_FSM_ERROR 3
`define DATA_WIDTH 32
