//
//------------------------------------------------------------------------------
//   Copyright 2018 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------------------------
//
//------------------------------------------------------------------------------
//   Copyright 2018 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------------------------
//----------------------------------------------------------------------
//   THIS IS AUTOMATICALLY GENERATED CODE
//   Generated by Mentor Graphics' Register Assistant UVM V4.6 (Build 8)
//   UVM Register Kit version 1.1
//----------------------------------------------------------------------
// Project         : PSS
// Unit            : pss_reg_pkg
// File            : pss_reg_pkg.sv
//----------------------------------------------------------------------
// Created by      : cgales
// Creation Date   : 2/11/16 12:55 PM
//----------------------------------------------------------------------
// Title           : PSS
//
// Description     :
//
//----------------------------------------------------------------------

//----------------------------------------------------------------------
// pss_reg_pkg
//----------------------------------------------------------------------
package pss_reg_pkg;

   import uvm_pkg::*;
   import spi_reg_pkg::*;
   import gpio_reg_pkg::*;

   `include "uvm_macros.svh"

   //--------------------------------------------------------------------
   // Class: sw_top_block
   //
   // Top block for the stopwatch design
   //--------------------------------------------------------------------

   class pss_reg_block extends uvm_reg_block;
      `uvm_object_utils(pss_reg_block)

      rand spi_reg_block spi_rb; // SPI register block
      rand gpio_reg_block gpio_rb; // GPIO register block

      uvm_reg_map pss_map; // PSS block map

      // Function: new
      //
      function new(string name = "pss_reg_block");
         super.new(name, build_coverage(UVM_CVR_ALL));
      endfunction

      // Function: build
      //
      virtual function void build();

         add_hdl_path("top.dut");

         spi_rb = spi_reg_block::type_id::create("spi_rb");
         spi_rb.configure(this);
         spi_rb.build();

         gpio_rb = gpio_reg_block::type_id::create("gpio_rb");
         gpio_rb.configure(this);
         gpio_rb.build();

         pss_map = create_map("pss_map", 'h0, 4, UVM_LITTLE_ENDIAN, 1);
         default_map = pss_map;

         pss_map.add_submap(spi_rb.spi_reg_block_map, 'h0);
         pss_map.add_submap(gpio_rb.gpio_reg_block_map, 'h0100);

         lock_model();
      endfunction

      // Function: sample
      //
      function void sample(uvm_reg_addr_t offset, bit is_read, uvm_reg_map  map);

      endfunction: sample

   endclass


endpackage
