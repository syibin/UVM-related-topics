//------------------------------------------------------------
//   Copyright 2010-2018 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------
package apb_slave_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

//import register_layering_pkg::*;

`include "apb_slave_seq_item.svh"
`include "apb_slave_agent_config.svh"
`include "apb_slave_driver.svh"
`include "apb_slave_monitor.svh"
`include "apb_slave_sequencer.svh"
`include "apb_listener.svh"
`include "apb_slave_agent.svh"

// Utility Sequences
`include "apb_slave_sequence.svh"

endpackage: apb_slave_agent_pkg
